##
## LEF for PtnCells ;
## created by Encounter v09.10-p004_1 on Thu Nov 21 10:50:50 2013
##

VERSION 5.5 ;

NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

UNITS
  DATABASE MICRONS 2000 ;
END UNITS

MACRO RegFile
  CLASS BLOCK ;
  SIZE 89.7700 BY 89.2600 ;
  FOREIGN RegFile 0.0000 0.0000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN addressA[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 32.7400 89.1900 32.8100 89.2600 ;
    END
  END addressA[4]
  PIN addressA[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 31.7900 89.1900 31.8600 89.2600 ;
    END
  END addressA[3]
  PIN addressA[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 30.8400 89.1900 30.9100 89.2600 ;
    END
  END addressA[2]
  PIN addressA[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 29.8900 89.1900 29.9600 89.2600 ;
    END
  END addressA[1]
  PIN addressA[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 28.9400 89.1900 29.0100 89.2600 ;
    END
  END addressA[0]
  PIN addressB[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 37.4900 89.1900 37.5600 89.2600 ;
    END
  END addressB[4]
  PIN addressB[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 36.5400 89.1900 36.6100 89.2600 ;
    END
  END addressB[3]
  PIN addressB[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 35.5900 89.1900 35.6600 89.2600 ;
    END
  END addressB[2]
  PIN addressB[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 34.6400 89.1900 34.7100 89.2600 ;
    END
  END addressB[1]
  PIN addressB[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 33.6900 89.1900 33.7600 89.2600 ;
    END
  END addressB[0]
  PIN dataIn[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 52.6900 89.1900 52.7600 89.2600 ;
    END
  END dataIn[15]
  PIN dataIn[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 51.7400 89.1900 51.8100 89.2600 ;
    END
  END dataIn[14]
  PIN dataIn[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 50.7900 89.1900 50.8600 89.2600 ;
    END
  END dataIn[13]
  PIN dataIn[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 49.8400 89.1900 49.9100 89.2600 ;
    END
  END dataIn[12]
  PIN dataIn[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 48.8900 89.1900 48.9600 89.2600 ;
    END
  END dataIn[11]
  PIN dataIn[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 47.9400 89.1900 48.0100 89.2600 ;
    END
  END dataIn[10]
  PIN dataIn[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 62.7600 0.0000 62.8300 0.0700 ;
    END
  END dataIn[9]
  PIN dataIn[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 46.0400 89.1900 46.1100 89.2600 ;
    END
  END dataIn[8]
  PIN dataIn[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 45.0900 89.1900 45.1600 89.2600 ;
    END
  END dataIn[7]
  PIN dataIn[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 44.1400 89.1900 44.2100 89.2600 ;
    END
  END dataIn[6]
  PIN dataIn[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 43.1900 89.1900 43.2600 89.2600 ;
    END
  END dataIn[5]
  PIN dataIn[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 42.2400 89.1900 42.3100 89.2600 ;
    END
  END dataIn[4]
  PIN dataIn[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 41.2900 89.1900 41.3600 89.2600 ;
    END
  END dataIn[3]
  PIN dataIn[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 40.3400 89.1900 40.4100 89.2600 ;
    END
  END dataIn[2]
  PIN dataIn[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 39.3900 89.1900 39.4600 89.2600 ;
    END
  END dataIn[1]
  PIN dataIn[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 38.4400 89.1900 38.5100 89.2600 ;
    END
  END dataIn[0]
  PIN addressIn[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 57.4400 89.1900 57.5100 89.2600 ;
    END
  END addressIn[4]
  PIN addressIn[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 56.4900 89.1900 56.5600 89.2600 ;
    END
  END addressIn[3]
  PIN addressIn[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 55.5400 89.1900 55.6100 89.2600 ;
    END
  END addressIn[2]
  PIN addressIn[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 54.5900 89.1900 54.6600 89.2600 ;
    END
  END addressIn[1]
  PIN addressIn[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 53.6400 89.1900 53.7100 89.2600 ;
    END
  END addressIn[0]
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 58.3900 89.1900 58.4600 89.2600 ;
    END
  END clk
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 59.3400 89.1900 59.4100 89.2600 ;
    END
  END reset
  PIN write
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 60.2900 89.1900 60.3600 89.2600 ;
    END
  END write
  PIN outA[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 43.7600 0.0000 43.8300 0.0700 ;
    END
  END outA[15]
  PIN outA[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 41.8600 0.0000 41.9300 0.0700 ;
    END
  END outA[14]
  PIN outA[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 39.9600 0.0000 40.0300 0.0700 ;
    END
  END outA[13]
  PIN outA[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 38.0600 0.0000 38.1300 0.0700 ;
    END
  END outA[12]
  PIN outA[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 36.1600 0.0000 36.2300 0.0700 ;
    END
  END outA[11]
  PIN outA[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 34.2600 0.0000 34.3300 0.0700 ;
    END
  END outA[10]
  PIN outA[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 32.3600 0.0000 32.4300 0.0700 ;
    END
  END outA[9]
  PIN outA[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 30.4600 0.0000 30.5300 0.0700 ;
    END
  END outA[8]
  PIN outA[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 28.5600 0.0000 28.6300 0.0700 ;
    END
  END outA[7]
  PIN outA[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 26.6600 0.0000 26.7300 0.0700 ;
    END
  END outA[6]
  PIN outA[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 24.7600 0.0000 24.8300 0.0700 ;
    END
  END outA[5]
  PIN outA[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 22.8600 0.0000 22.9300 0.0700 ;
    END
  END outA[4]
  PIN outA[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 20.9600 0.0000 21.0300 0.0700 ;
    END
  END outA[3]
  PIN outA[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 19.0600 0.0000 19.1300 0.0700 ;
    END
  END outA[2]
  PIN outA[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 17.1600 0.0000 17.2300 0.0700 ;
    END
  END outA[1]
  PIN outA[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 15.2600 0.0000 15.3300 0.0700 ;
    END
  END outA[0]
  PIN outB[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 74.1600 0.0000 74.2300 0.0700 ;
    END
  END outB[15]
  PIN outB[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 72.2600 0.0000 72.3300 0.0700 ;
    END
  END outB[14]
  PIN outB[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 70.3600 0.0000 70.4300 0.0700 ;
    END
  END outB[13]
  PIN outB[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 68.4600 0.0000 68.5300 0.0700 ;
    END
  END outB[12]
  PIN outB[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 66.5600 0.0000 66.6300 0.0700 ;
    END
  END outB[11]
  PIN outB[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 64.6600 0.0000 64.7300 0.0700 ;
    END
  END outB[10]
  PIN outB[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 48.5100 0.0000 48.5800 0.0700 ;
    END
  END outB[9]
  PIN outB[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 60.8600 0.0000 60.9300 0.0700 ;
    END
  END outB[8]
  PIN outB[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 58.9600 0.0000 59.0300 0.0700 ;
    END
  END outB[7]
  PIN outB[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 57.0600 0.0000 57.1300 0.0700 ;
    END
  END outB[6]
  PIN outB[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 55.1600 0.0000 55.2300 0.0700 ;
    END
  END outB[5]
  PIN outB[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 53.2600 0.0000 53.3300 0.0700 ;
    END
  END outB[4]
  PIN outB[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 51.3600 0.0000 51.4300 0.0700 ;
    END
  END outB[3]
  PIN outB[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 49.4600 0.0000 49.5300 0.0700 ;
    END
  END outB[2]
  PIN outB[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 47.5600 0.0000 47.6300 0.0700 ;
    END
  END outB[1]
  PIN outB[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 45.6600 0.0000 45.7300 0.0700 ;
    END
  END outB[0]
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal10 ;
        RECT 86.6900 88.4600 87.4900 89.2600 ;
    END
    PORT
      LAYER metal10 ;
        RECT 86.6900 0.0000 87.4900 0.8000 ;
    END
    PORT
      LAYER metal10 ;
        RECT 2.3800 88.4600 3.1800 89.2600 ;
    END
    PORT
      LAYER metal10 ;
        RECT 2.3800 0.0000 3.1800 0.8000 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal10 ;
        RECT 88.2900 88.4600 89.0900 89.2600 ;
    END
    PORT
      LAYER metal10 ;
        RECT 88.2900 0.0000 89.0900 0.8000 ;
    END
    PORT
      LAYER metal10 ;
        RECT 0.7800 88.4600 1.5800 89.2600 ;
    END
    PORT
      LAYER metal10 ;
        RECT 0.7800 0.0000 1.5800 0.8000 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.0000 0.0000 89.7700 89.2600 ;
    LAYER metal2 ;
      RECT 60.4300 89.1200 89.7700 89.2600 ;
      RECT 59.4800 89.1200 60.2200 89.2600 ;
      RECT 58.5300 89.1200 59.2700 89.2600 ;
      RECT 57.5800 89.1200 58.3200 89.2600 ;
      RECT 56.6300 89.1200 57.3700 89.2600 ;
      RECT 55.6800 89.1200 56.4200 89.2600 ;
      RECT 54.7300 89.1200 55.4700 89.2600 ;
      RECT 53.7800 89.1200 54.5200 89.2600 ;
      RECT 52.8300 89.1200 53.5700 89.2600 ;
      RECT 51.8800 89.1200 52.6200 89.2600 ;
      RECT 50.9300 89.1200 51.6700 89.2600 ;
      RECT 49.9800 89.1200 50.7200 89.2600 ;
      RECT 49.0300 89.1200 49.7700 89.2600 ;
      RECT 48.0800 89.1200 48.8200 89.2600 ;
      RECT 46.1800 89.1200 47.8700 89.2600 ;
      RECT 45.2300 89.1200 45.9700 89.2600 ;
      RECT 44.2800 89.1200 45.0200 89.2600 ;
      RECT 43.3300 89.1200 44.0700 89.2600 ;
      RECT 42.3800 89.1200 43.1200 89.2600 ;
      RECT 41.4300 89.1200 42.1700 89.2600 ;
      RECT 40.4800 89.1200 41.2200 89.2600 ;
      RECT 39.5300 89.1200 40.2700 89.2600 ;
      RECT 38.5800 89.1200 39.3200 89.2600 ;
      RECT 37.6300 89.1200 38.3700 89.2600 ;
      RECT 36.6800 89.1200 37.4200 89.2600 ;
      RECT 35.7300 89.1200 36.4700 89.2600 ;
      RECT 34.7800 89.1200 35.5200 89.2600 ;
      RECT 33.8300 89.1200 34.5700 89.2600 ;
      RECT 32.8800 89.1200 33.6200 89.2600 ;
      RECT 31.9300 89.1200 32.6700 89.2600 ;
      RECT 30.9800 89.1200 31.7200 89.2600 ;
      RECT 30.0300 89.1200 30.7700 89.2600 ;
      RECT 29.0800 89.1200 29.8200 89.2600 ;
      RECT 0.0000 89.1200 28.8700 89.2600 ;
      RECT 0.0000 0.1400 89.7700 89.1200 ;
      RECT 74.3000 0.0000 89.7700 0.1400 ;
      RECT 72.4000 0.0000 74.0900 0.1400 ;
      RECT 70.5000 0.0000 72.1900 0.1400 ;
      RECT 68.6000 0.0000 70.2900 0.1400 ;
      RECT 66.7000 0.0000 68.3900 0.1400 ;
      RECT 64.8000 0.0000 66.4900 0.1400 ;
      RECT 62.9000 0.0000 64.5900 0.1400 ;
      RECT 61.0000 0.0000 62.6900 0.1400 ;
      RECT 59.1000 0.0000 60.7900 0.1400 ;
      RECT 57.2000 0.0000 58.8900 0.1400 ;
      RECT 55.3000 0.0000 56.9900 0.1400 ;
      RECT 53.4000 0.0000 55.0900 0.1400 ;
      RECT 51.5000 0.0000 53.1900 0.1400 ;
      RECT 49.6000 0.0000 51.2900 0.1400 ;
      RECT 48.6500 0.0000 49.3900 0.1400 ;
      RECT 47.7000 0.0000 48.4400 0.1400 ;
      RECT 45.8000 0.0000 47.4900 0.1400 ;
      RECT 43.9000 0.0000 45.5900 0.1400 ;
      RECT 42.0000 0.0000 43.6900 0.1400 ;
      RECT 40.1000 0.0000 41.7900 0.1400 ;
      RECT 38.2000 0.0000 39.8900 0.1400 ;
      RECT 36.3000 0.0000 37.9900 0.1400 ;
      RECT 34.4000 0.0000 36.0900 0.1400 ;
      RECT 32.5000 0.0000 34.1900 0.1400 ;
      RECT 30.6000 0.0000 32.2900 0.1400 ;
      RECT 28.7000 0.0000 30.3900 0.1400 ;
      RECT 26.8000 0.0000 28.4900 0.1400 ;
      RECT 24.9000 0.0000 26.5900 0.1400 ;
      RECT 23.0000 0.0000 24.6900 0.1400 ;
      RECT 21.1000 0.0000 22.7900 0.1400 ;
      RECT 19.2000 0.0000 20.8900 0.1400 ;
      RECT 17.3000 0.0000 18.9900 0.1400 ;
      RECT 15.4000 0.0000 17.0900 0.1400 ;
      RECT 0.0000 0.0000 15.1900 0.1400 ;
    LAYER metal3 ;
      RECT 0.0000 0.0000 89.7700 89.2600 ;
    LAYER metal4 ;
      RECT 0.0000 0.0000 89.7700 89.2600 ;
    LAYER metal5 ;
      RECT 0.0000 0.0000 89.7700 89.2600 ;
    LAYER metal6 ;
      RECT 0.0000 0.0000 89.7700 89.2600 ;
    LAYER metal7 ;
      RECT 0.0000 0.0000 89.7700 89.2600 ;
    LAYER metal8 ;
      RECT 0.0000 0.0000 89.7700 89.2600 ;
    LAYER metal9 ;
      RECT 0.0000 0.0000 89.7700 89.2600 ;
    LAYER metal10 ;
      RECT 3.9800 87.6600 85.8900 89.2600 ;
      RECT 0.0000 1.6000 89.7700 87.6600 ;
      RECT 3.9800 0.0000 85.8900 1.6000 ;
  END
END RegFile

END LIBRARY
