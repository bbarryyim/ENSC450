
module SingleReg_30 ( data, clk, reset, write, dataOut );
  input [15:0] data;
  output [15:0] dataOut;
  input clk, reset, write;
  wire   n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n100, n101;

  DFFR_X1 \Reg_reg[15]  ( .D(n53), .CK(clk), .RN(n54), .Q(dataOut[15]), .QN(
        n70) );
  DFFR_X1 \Reg_reg[14]  ( .D(n55), .CK(clk), .RN(n54), .Q(dataOut[14]), .QN(
        n71) );
  DFFR_X1 \Reg_reg[13]  ( .D(n56), .CK(clk), .RN(n54), .Q(dataOut[13]), .QN(
        n72) );
  DFFR_X1 \Reg_reg[12]  ( .D(n57), .CK(clk), .RN(n54), .Q(dataOut[12]), .QN(
        n73) );
  DFFR_X1 \Reg_reg[11]  ( .D(n58), .CK(clk), .RN(n54), .Q(dataOut[11]), .QN(
        n74) );
  DFFR_X1 \Reg_reg[10]  ( .D(n59), .CK(clk), .RN(n54), .Q(dataOut[10]), .QN(
        n75) );
  DFFR_X1 \Reg_reg[9]  ( .D(n60), .CK(clk), .RN(n54), .Q(dataOut[9]), .QN(n76)
         );
  DFFR_X1 \Reg_reg[8]  ( .D(n61), .CK(clk), .RN(n54), .Q(dataOut[8]), .QN(n77)
         );
  DFFR_X1 \Reg_reg[7]  ( .D(n62), .CK(clk), .RN(n54), .Q(dataOut[7]), .QN(n78)
         );
  DFFR_X1 \Reg_reg[6]  ( .D(n63), .CK(clk), .RN(n54), .Q(dataOut[6]), .QN(n79)
         );
  DFFR_X1 \Reg_reg[5]  ( .D(n64), .CK(clk), .RN(n54), .Q(dataOut[5]), .QN(n80)
         );
  DFFR_X1 \Reg_reg[4]  ( .D(n65), .CK(clk), .RN(n54), .Q(dataOut[4]), .QN(n81)
         );
  DFFR_X1 \Reg_reg[3]  ( .D(n66), .CK(clk), .RN(n54), .Q(dataOut[3]), .QN(n82)
         );
  DFFR_X1 \Reg_reg[2]  ( .D(n67), .CK(clk), .RN(n54), .Q(dataOut[2]), .QN(n83)
         );
  DFFR_X1 \Reg_reg[1]  ( .D(n68), .CK(clk), .RN(n54), .Q(dataOut[1]), .QN(n84)
         );
  DFFR_X1 \Reg_reg[0]  ( .D(n69), .CK(clk), .RN(n54), .Q(dataOut[0]), .QN(n85)
         );
  OAI21_X1 U2 ( .B1(n50), .B2(n85), .A(n101), .ZN(n69) );
  NAND2_X1 U3 ( .A1(n52), .A2(data[0]), .ZN(n101) );
  OAI21_X1 U4 ( .B1(n50), .B2(n84), .A(n100), .ZN(n68) );
  NAND2_X1 U5 ( .A1(data[1]), .A2(n52), .ZN(n100) );
  OAI21_X1 U6 ( .B1(n50), .B2(n83), .A(n99), .ZN(n67) );
  NAND2_X1 U7 ( .A1(data[2]), .A2(n52), .ZN(n99) );
  OAI21_X1 U8 ( .B1(n50), .B2(n82), .A(n98), .ZN(n66) );
  NAND2_X1 U9 ( .A1(data[3]), .A2(n52), .ZN(n98) );
  OAI21_X1 U10 ( .B1(n50), .B2(n81), .A(n97), .ZN(n65) );
  NAND2_X1 U11 ( .A1(data[4]), .A2(n52), .ZN(n97) );
  OAI21_X1 U12 ( .B1(n50), .B2(n80), .A(n96), .ZN(n64) );
  NAND2_X1 U13 ( .A1(data[5]), .A2(n52), .ZN(n96) );
  OAI21_X1 U14 ( .B1(n50), .B2(n79), .A(n95), .ZN(n63) );
  NAND2_X1 U15 ( .A1(data[6]), .A2(n52), .ZN(n95) );
  OAI21_X1 U16 ( .B1(n51), .B2(n78), .A(n94), .ZN(n62) );
  NAND2_X1 U17 ( .A1(data[7]), .A2(n52), .ZN(n94) );
  OAI21_X1 U18 ( .B1(n51), .B2(n77), .A(n93), .ZN(n61) );
  NAND2_X1 U19 ( .A1(data[8]), .A2(n51), .ZN(n93) );
  OAI21_X1 U20 ( .B1(n51), .B2(n76), .A(n92), .ZN(n60) );
  NAND2_X1 U21 ( .A1(data[9]), .A2(n51), .ZN(n92) );
  OAI21_X1 U22 ( .B1(n50), .B2(n75), .A(n91), .ZN(n59) );
  NAND2_X1 U23 ( .A1(data[10]), .A2(n51), .ZN(n91) );
  OAI21_X1 U24 ( .B1(n51), .B2(n74), .A(n90), .ZN(n58) );
  NAND2_X1 U25 ( .A1(data[11]), .A2(n51), .ZN(n90) );
  OAI21_X1 U26 ( .B1(n50), .B2(n73), .A(n89), .ZN(n57) );
  NAND2_X1 U27 ( .A1(data[12]), .A2(n51), .ZN(n89) );
  OAI21_X1 U28 ( .B1(n50), .B2(n72), .A(n88), .ZN(n56) );
  NAND2_X1 U29 ( .A1(data[13]), .A2(n51), .ZN(n88) );
  OAI21_X1 U30 ( .B1(n50), .B2(n71), .A(n87), .ZN(n55) );
  NAND2_X1 U31 ( .A1(data[14]), .A2(n51), .ZN(n87) );
  INV_X1 U32 ( .A(reset), .ZN(n54) );
  OAI21_X1 U33 ( .B1(n50), .B2(n70), .A(n86), .ZN(n53) );
  NAND2_X1 U34 ( .A1(data[15]), .A2(n51), .ZN(n86) );
  CLKBUF_X3 U35 ( .A(write), .Z(n50) );
  CLKBUF_X3 U36 ( .A(write), .Z(n51) );
  CLKBUF_X3 U37 ( .A(write), .Z(n52) );
endmodule


module SingleReg_29 ( data, clk, reset, write, dataOut );
  input [15:0] data;
  output [15:0] dataOut;
  input clk, reset, write;
  wire   n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n100, n101;

  DFFR_X1 \Reg_reg[15]  ( .D(n53), .CK(clk), .RN(n54), .Q(dataOut[15]), .QN(
        n70) );
  DFFR_X1 \Reg_reg[14]  ( .D(n55), .CK(clk), .RN(n54), .Q(dataOut[14]), .QN(
        n71) );
  DFFR_X1 \Reg_reg[13]  ( .D(n56), .CK(clk), .RN(n54), .Q(dataOut[13]), .QN(
        n72) );
  DFFR_X1 \Reg_reg[12]  ( .D(n57), .CK(clk), .RN(n54), .Q(dataOut[12]), .QN(
        n73) );
  DFFR_X1 \Reg_reg[11]  ( .D(n58), .CK(clk), .RN(n54), .Q(dataOut[11]), .QN(
        n74) );
  DFFR_X1 \Reg_reg[10]  ( .D(n59), .CK(clk), .RN(n54), .Q(dataOut[10]), .QN(
        n75) );
  DFFR_X1 \Reg_reg[9]  ( .D(n60), .CK(clk), .RN(n54), .Q(dataOut[9]), .QN(n76)
         );
  DFFR_X1 \Reg_reg[8]  ( .D(n61), .CK(clk), .RN(n54), .Q(dataOut[8]), .QN(n77)
         );
  DFFR_X1 \Reg_reg[7]  ( .D(n62), .CK(clk), .RN(n54), .Q(dataOut[7]), .QN(n78)
         );
  DFFR_X1 \Reg_reg[6]  ( .D(n63), .CK(clk), .RN(n54), .Q(dataOut[6]), .QN(n79)
         );
  DFFR_X1 \Reg_reg[5]  ( .D(n64), .CK(clk), .RN(n54), .Q(dataOut[5]), .QN(n80)
         );
  DFFR_X1 \Reg_reg[4]  ( .D(n65), .CK(clk), .RN(n54), .Q(dataOut[4]), .QN(n81)
         );
  DFFR_X1 \Reg_reg[3]  ( .D(n66), .CK(clk), .RN(n54), .Q(dataOut[3]), .QN(n82)
         );
  DFFR_X1 \Reg_reg[2]  ( .D(n67), .CK(clk), .RN(n54), .Q(dataOut[2]), .QN(n83)
         );
  DFFR_X1 \Reg_reg[1]  ( .D(n68), .CK(clk), .RN(n54), .Q(dataOut[1]), .QN(n84)
         );
  DFFR_X1 \Reg_reg[0]  ( .D(n69), .CK(clk), .RN(n54), .Q(dataOut[0]), .QN(n85)
         );
  OAI21_X1 U2 ( .B1(n50), .B2(n85), .A(n101), .ZN(n69) );
  NAND2_X1 U3 ( .A1(n52), .A2(data[0]), .ZN(n101) );
  OAI21_X1 U4 ( .B1(n50), .B2(n84), .A(n100), .ZN(n68) );
  NAND2_X1 U5 ( .A1(data[1]), .A2(n52), .ZN(n100) );
  OAI21_X1 U6 ( .B1(n50), .B2(n83), .A(n99), .ZN(n67) );
  NAND2_X1 U7 ( .A1(data[2]), .A2(n52), .ZN(n99) );
  OAI21_X1 U8 ( .B1(n50), .B2(n82), .A(n98), .ZN(n66) );
  NAND2_X1 U9 ( .A1(data[3]), .A2(n52), .ZN(n98) );
  OAI21_X1 U10 ( .B1(n50), .B2(n81), .A(n97), .ZN(n65) );
  NAND2_X1 U11 ( .A1(data[4]), .A2(n52), .ZN(n97) );
  OAI21_X1 U12 ( .B1(n50), .B2(n80), .A(n96), .ZN(n64) );
  NAND2_X1 U13 ( .A1(data[5]), .A2(n52), .ZN(n96) );
  OAI21_X1 U14 ( .B1(n50), .B2(n79), .A(n95), .ZN(n63) );
  NAND2_X1 U15 ( .A1(data[6]), .A2(n52), .ZN(n95) );
  OAI21_X1 U16 ( .B1(n51), .B2(n78), .A(n94), .ZN(n62) );
  NAND2_X1 U17 ( .A1(data[7]), .A2(n52), .ZN(n94) );
  OAI21_X1 U18 ( .B1(n51), .B2(n77), .A(n93), .ZN(n61) );
  NAND2_X1 U19 ( .A1(data[8]), .A2(n51), .ZN(n93) );
  OAI21_X1 U20 ( .B1(n51), .B2(n76), .A(n92), .ZN(n60) );
  NAND2_X1 U21 ( .A1(data[9]), .A2(n51), .ZN(n92) );
  OAI21_X1 U22 ( .B1(n50), .B2(n75), .A(n91), .ZN(n59) );
  NAND2_X1 U23 ( .A1(data[10]), .A2(n51), .ZN(n91) );
  OAI21_X1 U24 ( .B1(n51), .B2(n74), .A(n90), .ZN(n58) );
  NAND2_X1 U25 ( .A1(data[11]), .A2(n51), .ZN(n90) );
  OAI21_X1 U26 ( .B1(n50), .B2(n73), .A(n89), .ZN(n57) );
  NAND2_X1 U27 ( .A1(data[12]), .A2(n51), .ZN(n89) );
  OAI21_X1 U28 ( .B1(n50), .B2(n72), .A(n88), .ZN(n56) );
  NAND2_X1 U29 ( .A1(data[13]), .A2(n51), .ZN(n88) );
  OAI21_X1 U30 ( .B1(n50), .B2(n71), .A(n87), .ZN(n55) );
  NAND2_X1 U31 ( .A1(data[14]), .A2(n51), .ZN(n87) );
  INV_X1 U32 ( .A(reset), .ZN(n54) );
  OAI21_X1 U33 ( .B1(n50), .B2(n70), .A(n86), .ZN(n53) );
  NAND2_X1 U34 ( .A1(data[15]), .A2(n51), .ZN(n86) );
  CLKBUF_X3 U35 ( .A(write), .Z(n50) );
  CLKBUF_X3 U36 ( .A(write), .Z(n51) );
  CLKBUF_X3 U37 ( .A(write), .Z(n52) );
endmodule


module SingleReg_28 ( data, clk, reset, write, dataOut );
  input [15:0] data;
  output [15:0] dataOut;
  input clk, reset, write;
  wire   n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n100, n101;

  DFFR_X1 \Reg_reg[15]  ( .D(n53), .CK(clk), .RN(n54), .Q(dataOut[15]), .QN(
        n70) );
  DFFR_X1 \Reg_reg[14]  ( .D(n55), .CK(clk), .RN(n54), .Q(dataOut[14]), .QN(
        n71) );
  DFFR_X1 \Reg_reg[13]  ( .D(n56), .CK(clk), .RN(n54), .Q(dataOut[13]), .QN(
        n72) );
  DFFR_X1 \Reg_reg[12]  ( .D(n57), .CK(clk), .RN(n54), .Q(dataOut[12]), .QN(
        n73) );
  DFFR_X1 \Reg_reg[11]  ( .D(n58), .CK(clk), .RN(n54), .Q(dataOut[11]), .QN(
        n74) );
  DFFR_X1 \Reg_reg[10]  ( .D(n59), .CK(clk), .RN(n54), .Q(dataOut[10]), .QN(
        n75) );
  DFFR_X1 \Reg_reg[9]  ( .D(n60), .CK(clk), .RN(n54), .Q(dataOut[9]), .QN(n76)
         );
  DFFR_X1 \Reg_reg[8]  ( .D(n61), .CK(clk), .RN(n54), .Q(dataOut[8]), .QN(n77)
         );
  DFFR_X1 \Reg_reg[7]  ( .D(n62), .CK(clk), .RN(n54), .Q(dataOut[7]), .QN(n78)
         );
  DFFR_X1 \Reg_reg[6]  ( .D(n63), .CK(clk), .RN(n54), .Q(dataOut[6]), .QN(n79)
         );
  DFFR_X1 \Reg_reg[5]  ( .D(n64), .CK(clk), .RN(n54), .Q(dataOut[5]), .QN(n80)
         );
  DFFR_X1 \Reg_reg[4]  ( .D(n65), .CK(clk), .RN(n54), .Q(dataOut[4]), .QN(n81)
         );
  DFFR_X1 \Reg_reg[3]  ( .D(n66), .CK(clk), .RN(n54), .Q(dataOut[3]), .QN(n82)
         );
  DFFR_X1 \Reg_reg[2]  ( .D(n67), .CK(clk), .RN(n54), .Q(dataOut[2]), .QN(n83)
         );
  DFFR_X1 \Reg_reg[1]  ( .D(n68), .CK(clk), .RN(n54), .Q(dataOut[1]), .QN(n84)
         );
  DFFR_X1 \Reg_reg[0]  ( .D(n69), .CK(clk), .RN(n54), .Q(dataOut[0]), .QN(n85)
         );
  OAI21_X1 U2 ( .B1(n50), .B2(n85), .A(n101), .ZN(n69) );
  NAND2_X1 U3 ( .A1(n52), .A2(data[0]), .ZN(n101) );
  OAI21_X1 U4 ( .B1(n50), .B2(n84), .A(n100), .ZN(n68) );
  NAND2_X1 U5 ( .A1(data[1]), .A2(n52), .ZN(n100) );
  OAI21_X1 U6 ( .B1(n50), .B2(n83), .A(n99), .ZN(n67) );
  NAND2_X1 U7 ( .A1(data[2]), .A2(n52), .ZN(n99) );
  OAI21_X1 U8 ( .B1(n50), .B2(n82), .A(n98), .ZN(n66) );
  NAND2_X1 U9 ( .A1(data[3]), .A2(n52), .ZN(n98) );
  OAI21_X1 U10 ( .B1(n50), .B2(n81), .A(n97), .ZN(n65) );
  NAND2_X1 U11 ( .A1(data[4]), .A2(n52), .ZN(n97) );
  OAI21_X1 U12 ( .B1(n50), .B2(n80), .A(n96), .ZN(n64) );
  NAND2_X1 U13 ( .A1(data[5]), .A2(n52), .ZN(n96) );
  OAI21_X1 U14 ( .B1(n50), .B2(n79), .A(n95), .ZN(n63) );
  NAND2_X1 U15 ( .A1(data[6]), .A2(n52), .ZN(n95) );
  OAI21_X1 U16 ( .B1(n51), .B2(n78), .A(n94), .ZN(n62) );
  NAND2_X1 U17 ( .A1(data[7]), .A2(n52), .ZN(n94) );
  OAI21_X1 U18 ( .B1(n51), .B2(n77), .A(n93), .ZN(n61) );
  NAND2_X1 U19 ( .A1(data[8]), .A2(n51), .ZN(n93) );
  OAI21_X1 U20 ( .B1(n51), .B2(n76), .A(n92), .ZN(n60) );
  NAND2_X1 U21 ( .A1(data[9]), .A2(n51), .ZN(n92) );
  OAI21_X1 U22 ( .B1(n50), .B2(n75), .A(n91), .ZN(n59) );
  NAND2_X1 U23 ( .A1(data[10]), .A2(n51), .ZN(n91) );
  OAI21_X1 U24 ( .B1(n51), .B2(n74), .A(n90), .ZN(n58) );
  NAND2_X1 U25 ( .A1(data[11]), .A2(n51), .ZN(n90) );
  OAI21_X1 U26 ( .B1(n50), .B2(n73), .A(n89), .ZN(n57) );
  NAND2_X1 U27 ( .A1(data[12]), .A2(n51), .ZN(n89) );
  OAI21_X1 U28 ( .B1(n50), .B2(n72), .A(n88), .ZN(n56) );
  NAND2_X1 U29 ( .A1(data[13]), .A2(n51), .ZN(n88) );
  OAI21_X1 U30 ( .B1(n50), .B2(n71), .A(n87), .ZN(n55) );
  NAND2_X1 U31 ( .A1(data[14]), .A2(n51), .ZN(n87) );
  INV_X1 U32 ( .A(reset), .ZN(n54) );
  OAI21_X1 U33 ( .B1(n50), .B2(n70), .A(n86), .ZN(n53) );
  NAND2_X1 U34 ( .A1(data[15]), .A2(n51), .ZN(n86) );
  CLKBUF_X3 U35 ( .A(write), .Z(n50) );
  CLKBUF_X3 U36 ( .A(write), .Z(n51) );
  CLKBUF_X3 U37 ( .A(write), .Z(n52) );
endmodule


module SingleReg_27 ( data, clk, reset, write, dataOut );
  input [15:0] data;
  output [15:0] dataOut;
  input clk, reset, write;
  wire   n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n100, n101;

  DFFR_X1 \Reg_reg[15]  ( .D(n53), .CK(clk), .RN(n54), .Q(dataOut[15]), .QN(
        n70) );
  DFFR_X1 \Reg_reg[14]  ( .D(n55), .CK(clk), .RN(n54), .Q(dataOut[14]), .QN(
        n71) );
  DFFR_X1 \Reg_reg[13]  ( .D(n56), .CK(clk), .RN(n54), .Q(dataOut[13]), .QN(
        n72) );
  DFFR_X1 \Reg_reg[12]  ( .D(n57), .CK(clk), .RN(n54), .Q(dataOut[12]), .QN(
        n73) );
  DFFR_X1 \Reg_reg[11]  ( .D(n58), .CK(clk), .RN(n54), .Q(dataOut[11]), .QN(
        n74) );
  DFFR_X1 \Reg_reg[10]  ( .D(n59), .CK(clk), .RN(n54), .Q(dataOut[10]), .QN(
        n75) );
  DFFR_X1 \Reg_reg[9]  ( .D(n60), .CK(clk), .RN(n54), .Q(dataOut[9]), .QN(n76)
         );
  DFFR_X1 \Reg_reg[8]  ( .D(n61), .CK(clk), .RN(n54), .Q(dataOut[8]), .QN(n77)
         );
  DFFR_X1 \Reg_reg[7]  ( .D(n62), .CK(clk), .RN(n54), .Q(dataOut[7]), .QN(n78)
         );
  DFFR_X1 \Reg_reg[6]  ( .D(n63), .CK(clk), .RN(n54), .Q(dataOut[6]), .QN(n79)
         );
  DFFR_X1 \Reg_reg[5]  ( .D(n64), .CK(clk), .RN(n54), .Q(dataOut[5]), .QN(n80)
         );
  DFFR_X1 \Reg_reg[4]  ( .D(n65), .CK(clk), .RN(n54), .Q(dataOut[4]), .QN(n81)
         );
  DFFR_X1 \Reg_reg[3]  ( .D(n66), .CK(clk), .RN(n54), .Q(dataOut[3]), .QN(n82)
         );
  DFFR_X1 \Reg_reg[2]  ( .D(n67), .CK(clk), .RN(n54), .Q(dataOut[2]), .QN(n83)
         );
  DFFR_X1 \Reg_reg[1]  ( .D(n68), .CK(clk), .RN(n54), .Q(dataOut[1]), .QN(n84)
         );
  DFFR_X1 \Reg_reg[0]  ( .D(n69), .CK(clk), .RN(n54), .Q(dataOut[0]), .QN(n85)
         );
  OAI21_X1 U2 ( .B1(n50), .B2(n85), .A(n101), .ZN(n69) );
  NAND2_X1 U3 ( .A1(n52), .A2(data[0]), .ZN(n101) );
  OAI21_X1 U4 ( .B1(n50), .B2(n84), .A(n100), .ZN(n68) );
  NAND2_X1 U5 ( .A1(data[1]), .A2(n52), .ZN(n100) );
  OAI21_X1 U6 ( .B1(n50), .B2(n83), .A(n99), .ZN(n67) );
  NAND2_X1 U7 ( .A1(data[2]), .A2(n52), .ZN(n99) );
  OAI21_X1 U8 ( .B1(n50), .B2(n82), .A(n98), .ZN(n66) );
  NAND2_X1 U9 ( .A1(data[3]), .A2(n52), .ZN(n98) );
  OAI21_X1 U10 ( .B1(n50), .B2(n81), .A(n97), .ZN(n65) );
  NAND2_X1 U11 ( .A1(data[4]), .A2(n52), .ZN(n97) );
  OAI21_X1 U12 ( .B1(n50), .B2(n80), .A(n96), .ZN(n64) );
  NAND2_X1 U13 ( .A1(data[5]), .A2(n52), .ZN(n96) );
  OAI21_X1 U14 ( .B1(n50), .B2(n79), .A(n95), .ZN(n63) );
  NAND2_X1 U15 ( .A1(data[6]), .A2(n52), .ZN(n95) );
  OAI21_X1 U16 ( .B1(n51), .B2(n78), .A(n94), .ZN(n62) );
  NAND2_X1 U17 ( .A1(data[7]), .A2(n52), .ZN(n94) );
  OAI21_X1 U18 ( .B1(n51), .B2(n77), .A(n93), .ZN(n61) );
  NAND2_X1 U19 ( .A1(data[8]), .A2(n51), .ZN(n93) );
  OAI21_X1 U20 ( .B1(n51), .B2(n76), .A(n92), .ZN(n60) );
  NAND2_X1 U21 ( .A1(data[9]), .A2(n51), .ZN(n92) );
  OAI21_X1 U22 ( .B1(n50), .B2(n75), .A(n91), .ZN(n59) );
  NAND2_X1 U23 ( .A1(data[10]), .A2(n51), .ZN(n91) );
  OAI21_X1 U24 ( .B1(n51), .B2(n74), .A(n90), .ZN(n58) );
  NAND2_X1 U25 ( .A1(data[11]), .A2(n51), .ZN(n90) );
  OAI21_X1 U26 ( .B1(n50), .B2(n73), .A(n89), .ZN(n57) );
  NAND2_X1 U27 ( .A1(data[12]), .A2(n51), .ZN(n89) );
  OAI21_X1 U28 ( .B1(n50), .B2(n72), .A(n88), .ZN(n56) );
  NAND2_X1 U29 ( .A1(data[13]), .A2(n51), .ZN(n88) );
  OAI21_X1 U30 ( .B1(n50), .B2(n71), .A(n87), .ZN(n55) );
  NAND2_X1 U31 ( .A1(data[14]), .A2(n51), .ZN(n87) );
  INV_X1 U32 ( .A(reset), .ZN(n54) );
  OAI21_X1 U33 ( .B1(n50), .B2(n70), .A(n86), .ZN(n53) );
  NAND2_X1 U34 ( .A1(data[15]), .A2(n51), .ZN(n86) );
  CLKBUF_X3 U35 ( .A(write), .Z(n50) );
  CLKBUF_X3 U36 ( .A(write), .Z(n51) );
  CLKBUF_X3 U37 ( .A(write), .Z(n52) );
endmodule


module SingleReg_26 ( data, clk, reset, write, dataOut );
  input [15:0] data;
  output [15:0] dataOut;
  input clk, reset, write;
  wire   n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n100, n101;

  DFFR_X1 \Reg_reg[15]  ( .D(n53), .CK(clk), .RN(n54), .Q(dataOut[15]), .QN(
        n70) );
  DFFR_X1 \Reg_reg[14]  ( .D(n55), .CK(clk), .RN(n54), .Q(dataOut[14]), .QN(
        n71) );
  DFFR_X1 \Reg_reg[13]  ( .D(n56), .CK(clk), .RN(n54), .Q(dataOut[13]), .QN(
        n72) );
  DFFR_X1 \Reg_reg[12]  ( .D(n57), .CK(clk), .RN(n54), .Q(dataOut[12]), .QN(
        n73) );
  DFFR_X1 \Reg_reg[11]  ( .D(n58), .CK(clk), .RN(n54), .Q(dataOut[11]), .QN(
        n74) );
  DFFR_X1 \Reg_reg[10]  ( .D(n59), .CK(clk), .RN(n54), .Q(dataOut[10]), .QN(
        n75) );
  DFFR_X1 \Reg_reg[9]  ( .D(n60), .CK(clk), .RN(n54), .Q(dataOut[9]), .QN(n76)
         );
  DFFR_X1 \Reg_reg[8]  ( .D(n61), .CK(clk), .RN(n54), .Q(dataOut[8]), .QN(n77)
         );
  DFFR_X1 \Reg_reg[7]  ( .D(n62), .CK(clk), .RN(n54), .Q(dataOut[7]), .QN(n78)
         );
  DFFR_X1 \Reg_reg[6]  ( .D(n63), .CK(clk), .RN(n54), .Q(dataOut[6]), .QN(n79)
         );
  DFFR_X1 \Reg_reg[5]  ( .D(n64), .CK(clk), .RN(n54), .Q(dataOut[5]), .QN(n80)
         );
  DFFR_X1 \Reg_reg[4]  ( .D(n65), .CK(clk), .RN(n54), .Q(dataOut[4]), .QN(n81)
         );
  DFFR_X1 \Reg_reg[3]  ( .D(n66), .CK(clk), .RN(n54), .Q(dataOut[3]), .QN(n82)
         );
  DFFR_X1 \Reg_reg[2]  ( .D(n67), .CK(clk), .RN(n54), .Q(dataOut[2]), .QN(n83)
         );
  DFFR_X1 \Reg_reg[1]  ( .D(n68), .CK(clk), .RN(n54), .Q(dataOut[1]), .QN(n84)
         );
  DFFR_X1 \Reg_reg[0]  ( .D(n69), .CK(clk), .RN(n54), .Q(dataOut[0]), .QN(n85)
         );
  OAI21_X1 U2 ( .B1(n50), .B2(n85), .A(n101), .ZN(n69) );
  NAND2_X1 U3 ( .A1(n52), .A2(data[0]), .ZN(n101) );
  OAI21_X1 U4 ( .B1(n50), .B2(n84), .A(n100), .ZN(n68) );
  NAND2_X1 U5 ( .A1(data[1]), .A2(n52), .ZN(n100) );
  OAI21_X1 U6 ( .B1(n50), .B2(n83), .A(n99), .ZN(n67) );
  NAND2_X1 U7 ( .A1(data[2]), .A2(n52), .ZN(n99) );
  OAI21_X1 U8 ( .B1(n50), .B2(n82), .A(n98), .ZN(n66) );
  NAND2_X1 U9 ( .A1(data[3]), .A2(n52), .ZN(n98) );
  OAI21_X1 U10 ( .B1(n50), .B2(n81), .A(n97), .ZN(n65) );
  NAND2_X1 U11 ( .A1(data[4]), .A2(n52), .ZN(n97) );
  OAI21_X1 U12 ( .B1(n50), .B2(n80), .A(n96), .ZN(n64) );
  NAND2_X1 U13 ( .A1(data[5]), .A2(n52), .ZN(n96) );
  OAI21_X1 U14 ( .B1(n50), .B2(n79), .A(n95), .ZN(n63) );
  NAND2_X1 U15 ( .A1(data[6]), .A2(n52), .ZN(n95) );
  OAI21_X1 U16 ( .B1(n51), .B2(n78), .A(n94), .ZN(n62) );
  NAND2_X1 U17 ( .A1(data[7]), .A2(n52), .ZN(n94) );
  OAI21_X1 U18 ( .B1(n51), .B2(n77), .A(n93), .ZN(n61) );
  NAND2_X1 U19 ( .A1(data[8]), .A2(n51), .ZN(n93) );
  OAI21_X1 U20 ( .B1(n51), .B2(n76), .A(n92), .ZN(n60) );
  NAND2_X1 U21 ( .A1(data[9]), .A2(n51), .ZN(n92) );
  OAI21_X1 U22 ( .B1(n50), .B2(n75), .A(n91), .ZN(n59) );
  NAND2_X1 U23 ( .A1(data[10]), .A2(n51), .ZN(n91) );
  OAI21_X1 U24 ( .B1(n51), .B2(n74), .A(n90), .ZN(n58) );
  NAND2_X1 U25 ( .A1(data[11]), .A2(n51), .ZN(n90) );
  OAI21_X1 U26 ( .B1(n50), .B2(n73), .A(n89), .ZN(n57) );
  NAND2_X1 U27 ( .A1(data[12]), .A2(n51), .ZN(n89) );
  OAI21_X1 U28 ( .B1(n50), .B2(n72), .A(n88), .ZN(n56) );
  NAND2_X1 U29 ( .A1(data[13]), .A2(n51), .ZN(n88) );
  OAI21_X1 U30 ( .B1(n50), .B2(n71), .A(n87), .ZN(n55) );
  NAND2_X1 U31 ( .A1(data[14]), .A2(n51), .ZN(n87) );
  INV_X1 U32 ( .A(reset), .ZN(n54) );
  OAI21_X1 U33 ( .B1(n50), .B2(n70), .A(n86), .ZN(n53) );
  NAND2_X1 U34 ( .A1(data[15]), .A2(n51), .ZN(n86) );
  CLKBUF_X3 U35 ( .A(write), .Z(n50) );
  CLKBUF_X3 U36 ( .A(write), .Z(n51) );
  CLKBUF_X3 U37 ( .A(write), .Z(n52) );
endmodule


module SingleReg_25 ( data, clk, reset, write, dataOut );
  input [15:0] data;
  output [15:0] dataOut;
  input clk, reset, write;
  wire   n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n100, n101;

  DFFR_X1 \Reg_reg[15]  ( .D(n53), .CK(clk), .RN(n54), .Q(dataOut[15]), .QN(
        n70) );
  DFFR_X1 \Reg_reg[14]  ( .D(n55), .CK(clk), .RN(n54), .Q(dataOut[14]), .QN(
        n71) );
  DFFR_X1 \Reg_reg[13]  ( .D(n56), .CK(clk), .RN(n54), .Q(dataOut[13]), .QN(
        n72) );
  DFFR_X1 \Reg_reg[12]  ( .D(n57), .CK(clk), .RN(n54), .Q(dataOut[12]), .QN(
        n73) );
  DFFR_X1 \Reg_reg[11]  ( .D(n58), .CK(clk), .RN(n54), .Q(dataOut[11]), .QN(
        n74) );
  DFFR_X1 \Reg_reg[10]  ( .D(n59), .CK(clk), .RN(n54), .Q(dataOut[10]), .QN(
        n75) );
  DFFR_X1 \Reg_reg[9]  ( .D(n60), .CK(clk), .RN(n54), .Q(dataOut[9]), .QN(n76)
         );
  DFFR_X1 \Reg_reg[8]  ( .D(n61), .CK(clk), .RN(n54), .Q(dataOut[8]), .QN(n77)
         );
  DFFR_X1 \Reg_reg[7]  ( .D(n62), .CK(clk), .RN(n54), .Q(dataOut[7]), .QN(n78)
         );
  DFFR_X1 \Reg_reg[6]  ( .D(n63), .CK(clk), .RN(n54), .Q(dataOut[6]), .QN(n79)
         );
  DFFR_X1 \Reg_reg[5]  ( .D(n64), .CK(clk), .RN(n54), .Q(dataOut[5]), .QN(n80)
         );
  DFFR_X1 \Reg_reg[4]  ( .D(n65), .CK(clk), .RN(n54), .Q(dataOut[4]), .QN(n81)
         );
  DFFR_X1 \Reg_reg[3]  ( .D(n66), .CK(clk), .RN(n54), .Q(dataOut[3]), .QN(n82)
         );
  DFFR_X1 \Reg_reg[2]  ( .D(n67), .CK(clk), .RN(n54), .Q(dataOut[2]), .QN(n83)
         );
  DFFR_X1 \Reg_reg[1]  ( .D(n68), .CK(clk), .RN(n54), .Q(dataOut[1]), .QN(n84)
         );
  DFFR_X1 \Reg_reg[0]  ( .D(n69), .CK(clk), .RN(n54), .Q(dataOut[0]), .QN(n85)
         );
  OAI21_X1 U2 ( .B1(n50), .B2(n85), .A(n101), .ZN(n69) );
  NAND2_X1 U3 ( .A1(n52), .A2(data[0]), .ZN(n101) );
  OAI21_X1 U4 ( .B1(n50), .B2(n84), .A(n100), .ZN(n68) );
  NAND2_X1 U5 ( .A1(data[1]), .A2(n52), .ZN(n100) );
  OAI21_X1 U6 ( .B1(n50), .B2(n83), .A(n99), .ZN(n67) );
  NAND2_X1 U7 ( .A1(data[2]), .A2(n52), .ZN(n99) );
  OAI21_X1 U8 ( .B1(n50), .B2(n82), .A(n98), .ZN(n66) );
  NAND2_X1 U9 ( .A1(data[3]), .A2(n52), .ZN(n98) );
  OAI21_X1 U10 ( .B1(n50), .B2(n81), .A(n97), .ZN(n65) );
  NAND2_X1 U11 ( .A1(data[4]), .A2(n52), .ZN(n97) );
  OAI21_X1 U12 ( .B1(n50), .B2(n80), .A(n96), .ZN(n64) );
  NAND2_X1 U13 ( .A1(data[5]), .A2(n52), .ZN(n96) );
  OAI21_X1 U14 ( .B1(n50), .B2(n79), .A(n95), .ZN(n63) );
  NAND2_X1 U15 ( .A1(data[6]), .A2(n52), .ZN(n95) );
  OAI21_X1 U16 ( .B1(n51), .B2(n78), .A(n94), .ZN(n62) );
  NAND2_X1 U17 ( .A1(data[7]), .A2(n52), .ZN(n94) );
  OAI21_X1 U18 ( .B1(n51), .B2(n77), .A(n93), .ZN(n61) );
  NAND2_X1 U19 ( .A1(data[8]), .A2(n51), .ZN(n93) );
  OAI21_X1 U20 ( .B1(n51), .B2(n76), .A(n92), .ZN(n60) );
  NAND2_X1 U21 ( .A1(data[9]), .A2(n51), .ZN(n92) );
  OAI21_X1 U22 ( .B1(n50), .B2(n75), .A(n91), .ZN(n59) );
  NAND2_X1 U23 ( .A1(data[10]), .A2(n51), .ZN(n91) );
  OAI21_X1 U24 ( .B1(n51), .B2(n74), .A(n90), .ZN(n58) );
  NAND2_X1 U25 ( .A1(data[11]), .A2(n51), .ZN(n90) );
  OAI21_X1 U26 ( .B1(n50), .B2(n73), .A(n89), .ZN(n57) );
  NAND2_X1 U27 ( .A1(data[12]), .A2(n51), .ZN(n89) );
  OAI21_X1 U28 ( .B1(n50), .B2(n72), .A(n88), .ZN(n56) );
  NAND2_X1 U29 ( .A1(data[13]), .A2(n51), .ZN(n88) );
  OAI21_X1 U30 ( .B1(n50), .B2(n71), .A(n87), .ZN(n55) );
  NAND2_X1 U31 ( .A1(data[14]), .A2(n51), .ZN(n87) );
  INV_X1 U32 ( .A(reset), .ZN(n54) );
  OAI21_X1 U33 ( .B1(n50), .B2(n70), .A(n86), .ZN(n53) );
  NAND2_X1 U34 ( .A1(data[15]), .A2(n51), .ZN(n86) );
  CLKBUF_X3 U35 ( .A(write), .Z(n50) );
  CLKBUF_X3 U36 ( .A(write), .Z(n51) );
  CLKBUF_X3 U37 ( .A(write), .Z(n52) );
endmodule


module SingleReg_24 ( data, clk, reset, write, dataOut );
  input [15:0] data;
  output [15:0] dataOut;
  input clk, reset, write;
  wire   n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n100, n101;

  DFFR_X1 \Reg_reg[15]  ( .D(n53), .CK(clk), .RN(n54), .Q(dataOut[15]), .QN(
        n70) );
  DFFR_X1 \Reg_reg[14]  ( .D(n55), .CK(clk), .RN(n54), .Q(dataOut[14]), .QN(
        n71) );
  DFFR_X1 \Reg_reg[13]  ( .D(n56), .CK(clk), .RN(n54), .Q(dataOut[13]), .QN(
        n72) );
  DFFR_X1 \Reg_reg[12]  ( .D(n57), .CK(clk), .RN(n54), .Q(dataOut[12]), .QN(
        n73) );
  DFFR_X1 \Reg_reg[11]  ( .D(n58), .CK(clk), .RN(n54), .Q(dataOut[11]), .QN(
        n74) );
  DFFR_X1 \Reg_reg[10]  ( .D(n59), .CK(clk), .RN(n54), .Q(dataOut[10]), .QN(
        n75) );
  DFFR_X1 \Reg_reg[9]  ( .D(n60), .CK(clk), .RN(n54), .Q(dataOut[9]), .QN(n76)
         );
  DFFR_X1 \Reg_reg[8]  ( .D(n61), .CK(clk), .RN(n54), .Q(dataOut[8]), .QN(n77)
         );
  DFFR_X1 \Reg_reg[7]  ( .D(n62), .CK(clk), .RN(n54), .Q(dataOut[7]), .QN(n78)
         );
  DFFR_X1 \Reg_reg[6]  ( .D(n63), .CK(clk), .RN(n54), .Q(dataOut[6]), .QN(n79)
         );
  DFFR_X1 \Reg_reg[5]  ( .D(n64), .CK(clk), .RN(n54), .Q(dataOut[5]), .QN(n80)
         );
  DFFR_X1 \Reg_reg[4]  ( .D(n65), .CK(clk), .RN(n54), .Q(dataOut[4]), .QN(n81)
         );
  DFFR_X1 \Reg_reg[3]  ( .D(n66), .CK(clk), .RN(n54), .Q(dataOut[3]), .QN(n82)
         );
  DFFR_X1 \Reg_reg[2]  ( .D(n67), .CK(clk), .RN(n54), .Q(dataOut[2]), .QN(n83)
         );
  DFFR_X1 \Reg_reg[1]  ( .D(n68), .CK(clk), .RN(n54), .Q(dataOut[1]), .QN(n84)
         );
  DFFR_X1 \Reg_reg[0]  ( .D(n69), .CK(clk), .RN(n54), .Q(dataOut[0]), .QN(n85)
         );
  OAI21_X1 U2 ( .B1(n50), .B2(n85), .A(n101), .ZN(n69) );
  NAND2_X1 U3 ( .A1(n52), .A2(data[0]), .ZN(n101) );
  OAI21_X1 U4 ( .B1(n50), .B2(n84), .A(n100), .ZN(n68) );
  NAND2_X1 U5 ( .A1(data[1]), .A2(n52), .ZN(n100) );
  OAI21_X1 U6 ( .B1(n50), .B2(n83), .A(n99), .ZN(n67) );
  NAND2_X1 U7 ( .A1(data[2]), .A2(n52), .ZN(n99) );
  OAI21_X1 U8 ( .B1(n50), .B2(n82), .A(n98), .ZN(n66) );
  NAND2_X1 U9 ( .A1(data[3]), .A2(n52), .ZN(n98) );
  OAI21_X1 U10 ( .B1(n50), .B2(n81), .A(n97), .ZN(n65) );
  NAND2_X1 U11 ( .A1(data[4]), .A2(n52), .ZN(n97) );
  OAI21_X1 U12 ( .B1(n50), .B2(n80), .A(n96), .ZN(n64) );
  NAND2_X1 U13 ( .A1(data[5]), .A2(n52), .ZN(n96) );
  OAI21_X1 U14 ( .B1(n50), .B2(n79), .A(n95), .ZN(n63) );
  NAND2_X1 U15 ( .A1(data[6]), .A2(n52), .ZN(n95) );
  OAI21_X1 U16 ( .B1(n51), .B2(n78), .A(n94), .ZN(n62) );
  NAND2_X1 U17 ( .A1(data[7]), .A2(n52), .ZN(n94) );
  OAI21_X1 U18 ( .B1(n51), .B2(n77), .A(n93), .ZN(n61) );
  NAND2_X1 U19 ( .A1(data[8]), .A2(n51), .ZN(n93) );
  OAI21_X1 U20 ( .B1(n51), .B2(n76), .A(n92), .ZN(n60) );
  NAND2_X1 U21 ( .A1(data[9]), .A2(n51), .ZN(n92) );
  OAI21_X1 U22 ( .B1(n50), .B2(n75), .A(n91), .ZN(n59) );
  NAND2_X1 U23 ( .A1(data[10]), .A2(n51), .ZN(n91) );
  OAI21_X1 U24 ( .B1(n51), .B2(n74), .A(n90), .ZN(n58) );
  NAND2_X1 U25 ( .A1(data[11]), .A2(n51), .ZN(n90) );
  OAI21_X1 U26 ( .B1(n50), .B2(n73), .A(n89), .ZN(n57) );
  NAND2_X1 U27 ( .A1(data[12]), .A2(n51), .ZN(n89) );
  OAI21_X1 U28 ( .B1(n50), .B2(n72), .A(n88), .ZN(n56) );
  NAND2_X1 U29 ( .A1(data[13]), .A2(n51), .ZN(n88) );
  OAI21_X1 U30 ( .B1(n50), .B2(n71), .A(n87), .ZN(n55) );
  NAND2_X1 U31 ( .A1(data[14]), .A2(n51), .ZN(n87) );
  INV_X1 U32 ( .A(reset), .ZN(n54) );
  OAI21_X1 U33 ( .B1(n50), .B2(n70), .A(n86), .ZN(n53) );
  NAND2_X1 U34 ( .A1(data[15]), .A2(n51), .ZN(n86) );
  CLKBUF_X3 U35 ( .A(write), .Z(n50) );
  CLKBUF_X3 U36 ( .A(write), .Z(n51) );
  CLKBUF_X3 U37 ( .A(write), .Z(n52) );
endmodule


module SingleReg_23 ( data, clk, reset, write, dataOut );
  input [15:0] data;
  output [15:0] dataOut;
  input clk, reset, write;
  wire   n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n100, n101;

  DFFR_X1 \Reg_reg[15]  ( .D(n53), .CK(clk), .RN(n54), .Q(dataOut[15]), .QN(
        n70) );
  DFFR_X1 \Reg_reg[14]  ( .D(n55), .CK(clk), .RN(n54), .Q(dataOut[14]), .QN(
        n71) );
  DFFR_X1 \Reg_reg[13]  ( .D(n56), .CK(clk), .RN(n54), .Q(dataOut[13]), .QN(
        n72) );
  DFFR_X1 \Reg_reg[12]  ( .D(n57), .CK(clk), .RN(n54), .Q(dataOut[12]), .QN(
        n73) );
  DFFR_X1 \Reg_reg[11]  ( .D(n58), .CK(clk), .RN(n54), .Q(dataOut[11]), .QN(
        n74) );
  DFFR_X1 \Reg_reg[10]  ( .D(n59), .CK(clk), .RN(n54), .Q(dataOut[10]), .QN(
        n75) );
  DFFR_X1 \Reg_reg[9]  ( .D(n60), .CK(clk), .RN(n54), .Q(dataOut[9]), .QN(n76)
         );
  DFFR_X1 \Reg_reg[8]  ( .D(n61), .CK(clk), .RN(n54), .Q(dataOut[8]), .QN(n77)
         );
  DFFR_X1 \Reg_reg[7]  ( .D(n62), .CK(clk), .RN(n54), .Q(dataOut[7]), .QN(n78)
         );
  DFFR_X1 \Reg_reg[6]  ( .D(n63), .CK(clk), .RN(n54), .Q(dataOut[6]), .QN(n79)
         );
  DFFR_X1 \Reg_reg[5]  ( .D(n64), .CK(clk), .RN(n54), .Q(dataOut[5]), .QN(n80)
         );
  DFFR_X1 \Reg_reg[4]  ( .D(n65), .CK(clk), .RN(n54), .Q(dataOut[4]), .QN(n81)
         );
  DFFR_X1 \Reg_reg[3]  ( .D(n66), .CK(clk), .RN(n54), .Q(dataOut[3]), .QN(n82)
         );
  DFFR_X1 \Reg_reg[2]  ( .D(n67), .CK(clk), .RN(n54), .Q(dataOut[2]), .QN(n83)
         );
  DFFR_X1 \Reg_reg[1]  ( .D(n68), .CK(clk), .RN(n54), .Q(dataOut[1]), .QN(n84)
         );
  DFFR_X1 \Reg_reg[0]  ( .D(n69), .CK(clk), .RN(n54), .Q(dataOut[0]), .QN(n85)
         );
  OAI21_X1 U2 ( .B1(n50), .B2(n85), .A(n101), .ZN(n69) );
  NAND2_X1 U3 ( .A1(n52), .A2(data[0]), .ZN(n101) );
  OAI21_X1 U4 ( .B1(n50), .B2(n84), .A(n100), .ZN(n68) );
  NAND2_X1 U5 ( .A1(data[1]), .A2(n52), .ZN(n100) );
  OAI21_X1 U6 ( .B1(n50), .B2(n83), .A(n99), .ZN(n67) );
  NAND2_X1 U7 ( .A1(data[2]), .A2(n52), .ZN(n99) );
  OAI21_X1 U8 ( .B1(n50), .B2(n82), .A(n98), .ZN(n66) );
  NAND2_X1 U9 ( .A1(data[3]), .A2(n52), .ZN(n98) );
  OAI21_X1 U10 ( .B1(n50), .B2(n81), .A(n97), .ZN(n65) );
  NAND2_X1 U11 ( .A1(data[4]), .A2(n52), .ZN(n97) );
  OAI21_X1 U12 ( .B1(n50), .B2(n80), .A(n96), .ZN(n64) );
  NAND2_X1 U13 ( .A1(data[5]), .A2(n52), .ZN(n96) );
  OAI21_X1 U14 ( .B1(n50), .B2(n79), .A(n95), .ZN(n63) );
  NAND2_X1 U15 ( .A1(data[6]), .A2(n52), .ZN(n95) );
  OAI21_X1 U16 ( .B1(n51), .B2(n78), .A(n94), .ZN(n62) );
  NAND2_X1 U17 ( .A1(data[7]), .A2(n52), .ZN(n94) );
  OAI21_X1 U18 ( .B1(n51), .B2(n77), .A(n93), .ZN(n61) );
  NAND2_X1 U19 ( .A1(data[8]), .A2(n51), .ZN(n93) );
  OAI21_X1 U20 ( .B1(n51), .B2(n76), .A(n92), .ZN(n60) );
  NAND2_X1 U21 ( .A1(data[9]), .A2(n51), .ZN(n92) );
  OAI21_X1 U22 ( .B1(n50), .B2(n75), .A(n91), .ZN(n59) );
  NAND2_X1 U23 ( .A1(data[10]), .A2(n51), .ZN(n91) );
  OAI21_X1 U24 ( .B1(n51), .B2(n74), .A(n90), .ZN(n58) );
  NAND2_X1 U25 ( .A1(data[11]), .A2(n51), .ZN(n90) );
  OAI21_X1 U26 ( .B1(n50), .B2(n73), .A(n89), .ZN(n57) );
  NAND2_X1 U27 ( .A1(data[12]), .A2(n51), .ZN(n89) );
  OAI21_X1 U28 ( .B1(n50), .B2(n72), .A(n88), .ZN(n56) );
  NAND2_X1 U29 ( .A1(data[13]), .A2(n51), .ZN(n88) );
  OAI21_X1 U30 ( .B1(n50), .B2(n71), .A(n87), .ZN(n55) );
  NAND2_X1 U31 ( .A1(data[14]), .A2(n51), .ZN(n87) );
  INV_X1 U32 ( .A(reset), .ZN(n54) );
  OAI21_X1 U33 ( .B1(n50), .B2(n70), .A(n86), .ZN(n53) );
  NAND2_X1 U34 ( .A1(data[15]), .A2(n51), .ZN(n86) );
  CLKBUF_X3 U35 ( .A(write), .Z(n50) );
  CLKBUF_X3 U36 ( .A(write), .Z(n51) );
  CLKBUF_X3 U37 ( .A(write), .Z(n52) );
endmodule


module SingleReg_22 ( data, clk, reset, write, dataOut );
  input [15:0] data;
  output [15:0] dataOut;
  input clk, reset, write;
  wire   n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n100, n101;

  DFFR_X1 \Reg_reg[15]  ( .D(n53), .CK(clk), .RN(n54), .Q(dataOut[15]), .QN(
        n70) );
  DFFR_X1 \Reg_reg[14]  ( .D(n55), .CK(clk), .RN(n54), .Q(dataOut[14]), .QN(
        n71) );
  DFFR_X1 \Reg_reg[13]  ( .D(n56), .CK(clk), .RN(n54), .Q(dataOut[13]), .QN(
        n72) );
  DFFR_X1 \Reg_reg[12]  ( .D(n57), .CK(clk), .RN(n54), .Q(dataOut[12]), .QN(
        n73) );
  DFFR_X1 \Reg_reg[11]  ( .D(n58), .CK(clk), .RN(n54), .Q(dataOut[11]), .QN(
        n74) );
  DFFR_X1 \Reg_reg[10]  ( .D(n59), .CK(clk), .RN(n54), .Q(dataOut[10]), .QN(
        n75) );
  DFFR_X1 \Reg_reg[9]  ( .D(n60), .CK(clk), .RN(n54), .Q(dataOut[9]), .QN(n76)
         );
  DFFR_X1 \Reg_reg[8]  ( .D(n61), .CK(clk), .RN(n54), .Q(dataOut[8]), .QN(n77)
         );
  DFFR_X1 \Reg_reg[7]  ( .D(n62), .CK(clk), .RN(n54), .Q(dataOut[7]), .QN(n78)
         );
  DFFR_X1 \Reg_reg[6]  ( .D(n63), .CK(clk), .RN(n54), .Q(dataOut[6]), .QN(n79)
         );
  DFFR_X1 \Reg_reg[5]  ( .D(n64), .CK(clk), .RN(n54), .Q(dataOut[5]), .QN(n80)
         );
  DFFR_X1 \Reg_reg[4]  ( .D(n65), .CK(clk), .RN(n54), .Q(dataOut[4]), .QN(n81)
         );
  DFFR_X1 \Reg_reg[3]  ( .D(n66), .CK(clk), .RN(n54), .Q(dataOut[3]), .QN(n82)
         );
  DFFR_X1 \Reg_reg[2]  ( .D(n67), .CK(clk), .RN(n54), .Q(dataOut[2]), .QN(n83)
         );
  DFFR_X1 \Reg_reg[1]  ( .D(n68), .CK(clk), .RN(n54), .Q(dataOut[1]), .QN(n84)
         );
  DFFR_X1 \Reg_reg[0]  ( .D(n69), .CK(clk), .RN(n54), .Q(dataOut[0]), .QN(n85)
         );
  OAI21_X1 U2 ( .B1(n50), .B2(n85), .A(n101), .ZN(n69) );
  NAND2_X1 U3 ( .A1(n52), .A2(data[0]), .ZN(n101) );
  OAI21_X1 U4 ( .B1(n50), .B2(n84), .A(n100), .ZN(n68) );
  NAND2_X1 U5 ( .A1(data[1]), .A2(n52), .ZN(n100) );
  OAI21_X1 U6 ( .B1(n50), .B2(n83), .A(n99), .ZN(n67) );
  NAND2_X1 U7 ( .A1(data[2]), .A2(n52), .ZN(n99) );
  OAI21_X1 U8 ( .B1(n50), .B2(n82), .A(n98), .ZN(n66) );
  NAND2_X1 U9 ( .A1(data[3]), .A2(n52), .ZN(n98) );
  OAI21_X1 U10 ( .B1(n50), .B2(n81), .A(n97), .ZN(n65) );
  NAND2_X1 U11 ( .A1(data[4]), .A2(n52), .ZN(n97) );
  OAI21_X1 U12 ( .B1(n50), .B2(n80), .A(n96), .ZN(n64) );
  NAND2_X1 U13 ( .A1(data[5]), .A2(n52), .ZN(n96) );
  OAI21_X1 U14 ( .B1(n50), .B2(n79), .A(n95), .ZN(n63) );
  NAND2_X1 U15 ( .A1(data[6]), .A2(n52), .ZN(n95) );
  OAI21_X1 U16 ( .B1(n51), .B2(n78), .A(n94), .ZN(n62) );
  NAND2_X1 U17 ( .A1(data[7]), .A2(n52), .ZN(n94) );
  OAI21_X1 U18 ( .B1(n51), .B2(n77), .A(n93), .ZN(n61) );
  NAND2_X1 U19 ( .A1(data[8]), .A2(n51), .ZN(n93) );
  OAI21_X1 U20 ( .B1(n51), .B2(n76), .A(n92), .ZN(n60) );
  NAND2_X1 U21 ( .A1(data[9]), .A2(n51), .ZN(n92) );
  OAI21_X1 U22 ( .B1(n50), .B2(n75), .A(n91), .ZN(n59) );
  NAND2_X1 U23 ( .A1(data[10]), .A2(n51), .ZN(n91) );
  OAI21_X1 U24 ( .B1(n51), .B2(n74), .A(n90), .ZN(n58) );
  NAND2_X1 U25 ( .A1(data[11]), .A2(n51), .ZN(n90) );
  OAI21_X1 U26 ( .B1(n50), .B2(n73), .A(n89), .ZN(n57) );
  NAND2_X1 U27 ( .A1(data[12]), .A2(n51), .ZN(n89) );
  OAI21_X1 U28 ( .B1(n50), .B2(n72), .A(n88), .ZN(n56) );
  NAND2_X1 U29 ( .A1(data[13]), .A2(n51), .ZN(n88) );
  OAI21_X1 U30 ( .B1(n50), .B2(n71), .A(n87), .ZN(n55) );
  NAND2_X1 U31 ( .A1(data[14]), .A2(n51), .ZN(n87) );
  INV_X1 U32 ( .A(reset), .ZN(n54) );
  OAI21_X1 U33 ( .B1(n50), .B2(n70), .A(n86), .ZN(n53) );
  NAND2_X1 U34 ( .A1(data[15]), .A2(n51), .ZN(n86) );
  CLKBUF_X3 U35 ( .A(write), .Z(n50) );
  CLKBUF_X3 U36 ( .A(write), .Z(n51) );
  CLKBUF_X3 U37 ( .A(write), .Z(n52) );
endmodule


module SingleReg_21 ( data, clk, reset, write, dataOut );
  input [15:0] data;
  output [15:0] dataOut;
  input clk, reset, write;
  wire   n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n100, n101;

  DFFR_X1 \Reg_reg[15]  ( .D(n53), .CK(clk), .RN(n54), .Q(dataOut[15]), .QN(
        n70) );
  DFFR_X1 \Reg_reg[14]  ( .D(n55), .CK(clk), .RN(n54), .Q(dataOut[14]), .QN(
        n71) );
  DFFR_X1 \Reg_reg[13]  ( .D(n56), .CK(clk), .RN(n54), .Q(dataOut[13]), .QN(
        n72) );
  DFFR_X1 \Reg_reg[12]  ( .D(n57), .CK(clk), .RN(n54), .Q(dataOut[12]), .QN(
        n73) );
  DFFR_X1 \Reg_reg[11]  ( .D(n58), .CK(clk), .RN(n54), .Q(dataOut[11]), .QN(
        n74) );
  DFFR_X1 \Reg_reg[10]  ( .D(n59), .CK(clk), .RN(n54), .Q(dataOut[10]), .QN(
        n75) );
  DFFR_X1 \Reg_reg[9]  ( .D(n60), .CK(clk), .RN(n54), .Q(dataOut[9]), .QN(n76)
         );
  DFFR_X1 \Reg_reg[8]  ( .D(n61), .CK(clk), .RN(n54), .Q(dataOut[8]), .QN(n77)
         );
  DFFR_X1 \Reg_reg[7]  ( .D(n62), .CK(clk), .RN(n54), .Q(dataOut[7]), .QN(n78)
         );
  DFFR_X1 \Reg_reg[6]  ( .D(n63), .CK(clk), .RN(n54), .Q(dataOut[6]), .QN(n79)
         );
  DFFR_X1 \Reg_reg[5]  ( .D(n64), .CK(clk), .RN(n54), .Q(dataOut[5]), .QN(n80)
         );
  DFFR_X1 \Reg_reg[4]  ( .D(n65), .CK(clk), .RN(n54), .Q(dataOut[4]), .QN(n81)
         );
  DFFR_X1 \Reg_reg[3]  ( .D(n66), .CK(clk), .RN(n54), .Q(dataOut[3]), .QN(n82)
         );
  DFFR_X1 \Reg_reg[2]  ( .D(n67), .CK(clk), .RN(n54), .Q(dataOut[2]), .QN(n83)
         );
  DFFR_X1 \Reg_reg[1]  ( .D(n68), .CK(clk), .RN(n54), .Q(dataOut[1]), .QN(n84)
         );
  DFFR_X1 \Reg_reg[0]  ( .D(n69), .CK(clk), .RN(n54), .Q(dataOut[0]), .QN(n85)
         );
  OAI21_X1 U2 ( .B1(n50), .B2(n85), .A(n101), .ZN(n69) );
  NAND2_X1 U3 ( .A1(n52), .A2(data[0]), .ZN(n101) );
  OAI21_X1 U4 ( .B1(n50), .B2(n84), .A(n100), .ZN(n68) );
  NAND2_X1 U5 ( .A1(data[1]), .A2(n52), .ZN(n100) );
  OAI21_X1 U6 ( .B1(n50), .B2(n83), .A(n99), .ZN(n67) );
  NAND2_X1 U7 ( .A1(data[2]), .A2(n52), .ZN(n99) );
  OAI21_X1 U8 ( .B1(n50), .B2(n82), .A(n98), .ZN(n66) );
  NAND2_X1 U9 ( .A1(data[3]), .A2(n52), .ZN(n98) );
  OAI21_X1 U10 ( .B1(n50), .B2(n81), .A(n97), .ZN(n65) );
  NAND2_X1 U11 ( .A1(data[4]), .A2(n52), .ZN(n97) );
  OAI21_X1 U12 ( .B1(n50), .B2(n80), .A(n96), .ZN(n64) );
  NAND2_X1 U13 ( .A1(data[5]), .A2(n52), .ZN(n96) );
  OAI21_X1 U14 ( .B1(n50), .B2(n79), .A(n95), .ZN(n63) );
  NAND2_X1 U15 ( .A1(data[6]), .A2(n52), .ZN(n95) );
  OAI21_X1 U16 ( .B1(n51), .B2(n78), .A(n94), .ZN(n62) );
  NAND2_X1 U17 ( .A1(data[7]), .A2(n52), .ZN(n94) );
  OAI21_X1 U18 ( .B1(n51), .B2(n77), .A(n93), .ZN(n61) );
  NAND2_X1 U19 ( .A1(data[8]), .A2(n51), .ZN(n93) );
  OAI21_X1 U20 ( .B1(n51), .B2(n76), .A(n92), .ZN(n60) );
  NAND2_X1 U21 ( .A1(data[9]), .A2(n51), .ZN(n92) );
  OAI21_X1 U22 ( .B1(n50), .B2(n75), .A(n91), .ZN(n59) );
  NAND2_X1 U23 ( .A1(data[10]), .A2(n51), .ZN(n91) );
  OAI21_X1 U24 ( .B1(n51), .B2(n74), .A(n90), .ZN(n58) );
  NAND2_X1 U25 ( .A1(data[11]), .A2(n51), .ZN(n90) );
  OAI21_X1 U26 ( .B1(n50), .B2(n73), .A(n89), .ZN(n57) );
  NAND2_X1 U27 ( .A1(data[12]), .A2(n51), .ZN(n89) );
  OAI21_X1 U28 ( .B1(n50), .B2(n72), .A(n88), .ZN(n56) );
  NAND2_X1 U29 ( .A1(data[13]), .A2(n51), .ZN(n88) );
  OAI21_X1 U30 ( .B1(n50), .B2(n71), .A(n87), .ZN(n55) );
  NAND2_X1 U31 ( .A1(data[14]), .A2(n51), .ZN(n87) );
  INV_X1 U32 ( .A(reset), .ZN(n54) );
  OAI21_X1 U33 ( .B1(n50), .B2(n70), .A(n86), .ZN(n53) );
  NAND2_X1 U34 ( .A1(data[15]), .A2(n51), .ZN(n86) );
  CLKBUF_X3 U35 ( .A(write), .Z(n50) );
  CLKBUF_X3 U36 ( .A(write), .Z(n51) );
  CLKBUF_X3 U37 ( .A(write), .Z(n52) );
endmodule


module SingleReg_20 ( data, clk, reset, write, dataOut );
  input [15:0] data;
  output [15:0] dataOut;
  input clk, reset, write;
  wire   n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n100, n101;

  DFFR_X1 \Reg_reg[15]  ( .D(n53), .CK(clk), .RN(n54), .Q(dataOut[15]), .QN(
        n70) );
  DFFR_X1 \Reg_reg[14]  ( .D(n55), .CK(clk), .RN(n54), .Q(dataOut[14]), .QN(
        n71) );
  DFFR_X1 \Reg_reg[13]  ( .D(n56), .CK(clk), .RN(n54), .Q(dataOut[13]), .QN(
        n72) );
  DFFR_X1 \Reg_reg[12]  ( .D(n57), .CK(clk), .RN(n54), .Q(dataOut[12]), .QN(
        n73) );
  DFFR_X1 \Reg_reg[11]  ( .D(n58), .CK(clk), .RN(n54), .Q(dataOut[11]), .QN(
        n74) );
  DFFR_X1 \Reg_reg[10]  ( .D(n59), .CK(clk), .RN(n54), .Q(dataOut[10]), .QN(
        n75) );
  DFFR_X1 \Reg_reg[9]  ( .D(n60), .CK(clk), .RN(n54), .Q(dataOut[9]), .QN(n76)
         );
  DFFR_X1 \Reg_reg[8]  ( .D(n61), .CK(clk), .RN(n54), .Q(dataOut[8]), .QN(n77)
         );
  DFFR_X1 \Reg_reg[7]  ( .D(n62), .CK(clk), .RN(n54), .Q(dataOut[7]), .QN(n78)
         );
  DFFR_X1 \Reg_reg[6]  ( .D(n63), .CK(clk), .RN(n54), .Q(dataOut[6]), .QN(n79)
         );
  DFFR_X1 \Reg_reg[5]  ( .D(n64), .CK(clk), .RN(n54), .Q(dataOut[5]), .QN(n80)
         );
  DFFR_X1 \Reg_reg[4]  ( .D(n65), .CK(clk), .RN(n54), .Q(dataOut[4]), .QN(n81)
         );
  DFFR_X1 \Reg_reg[3]  ( .D(n66), .CK(clk), .RN(n54), .Q(dataOut[3]), .QN(n82)
         );
  DFFR_X1 \Reg_reg[2]  ( .D(n67), .CK(clk), .RN(n54), .Q(dataOut[2]), .QN(n83)
         );
  DFFR_X1 \Reg_reg[1]  ( .D(n68), .CK(clk), .RN(n54), .Q(dataOut[1]), .QN(n84)
         );
  DFFR_X1 \Reg_reg[0]  ( .D(n69), .CK(clk), .RN(n54), .Q(dataOut[0]), .QN(n85)
         );
  OAI21_X1 U2 ( .B1(n50), .B2(n85), .A(n101), .ZN(n69) );
  NAND2_X1 U3 ( .A1(n52), .A2(data[0]), .ZN(n101) );
  OAI21_X1 U4 ( .B1(n50), .B2(n84), .A(n100), .ZN(n68) );
  NAND2_X1 U5 ( .A1(data[1]), .A2(n52), .ZN(n100) );
  OAI21_X1 U6 ( .B1(n50), .B2(n83), .A(n99), .ZN(n67) );
  NAND2_X1 U7 ( .A1(data[2]), .A2(n52), .ZN(n99) );
  OAI21_X1 U8 ( .B1(n50), .B2(n82), .A(n98), .ZN(n66) );
  NAND2_X1 U9 ( .A1(data[3]), .A2(n52), .ZN(n98) );
  OAI21_X1 U10 ( .B1(n50), .B2(n81), .A(n97), .ZN(n65) );
  NAND2_X1 U11 ( .A1(data[4]), .A2(n52), .ZN(n97) );
  OAI21_X1 U12 ( .B1(n50), .B2(n80), .A(n96), .ZN(n64) );
  NAND2_X1 U13 ( .A1(data[5]), .A2(n52), .ZN(n96) );
  OAI21_X1 U14 ( .B1(n50), .B2(n79), .A(n95), .ZN(n63) );
  NAND2_X1 U15 ( .A1(data[6]), .A2(n52), .ZN(n95) );
  OAI21_X1 U16 ( .B1(n51), .B2(n78), .A(n94), .ZN(n62) );
  NAND2_X1 U17 ( .A1(data[7]), .A2(n52), .ZN(n94) );
  OAI21_X1 U18 ( .B1(n51), .B2(n77), .A(n93), .ZN(n61) );
  NAND2_X1 U19 ( .A1(data[8]), .A2(n51), .ZN(n93) );
  OAI21_X1 U20 ( .B1(n51), .B2(n76), .A(n92), .ZN(n60) );
  NAND2_X1 U21 ( .A1(data[9]), .A2(n51), .ZN(n92) );
  OAI21_X1 U22 ( .B1(n50), .B2(n75), .A(n91), .ZN(n59) );
  NAND2_X1 U23 ( .A1(data[10]), .A2(n51), .ZN(n91) );
  OAI21_X1 U24 ( .B1(n51), .B2(n74), .A(n90), .ZN(n58) );
  NAND2_X1 U25 ( .A1(data[11]), .A2(n51), .ZN(n90) );
  OAI21_X1 U26 ( .B1(n50), .B2(n73), .A(n89), .ZN(n57) );
  NAND2_X1 U27 ( .A1(data[12]), .A2(n51), .ZN(n89) );
  OAI21_X1 U28 ( .B1(n50), .B2(n72), .A(n88), .ZN(n56) );
  NAND2_X1 U29 ( .A1(data[13]), .A2(n51), .ZN(n88) );
  OAI21_X1 U30 ( .B1(n50), .B2(n71), .A(n87), .ZN(n55) );
  NAND2_X1 U31 ( .A1(data[14]), .A2(n51), .ZN(n87) );
  INV_X1 U32 ( .A(reset), .ZN(n54) );
  OAI21_X1 U33 ( .B1(n50), .B2(n70), .A(n86), .ZN(n53) );
  NAND2_X1 U34 ( .A1(data[15]), .A2(n51), .ZN(n86) );
  CLKBUF_X3 U35 ( .A(write), .Z(n50) );
  CLKBUF_X3 U36 ( .A(write), .Z(n51) );
  CLKBUF_X3 U37 ( .A(write), .Z(n52) );
endmodule


module SingleReg_19 ( data, clk, reset, write, dataOut );
  input [15:0] data;
  output [15:0] dataOut;
  input clk, reset, write;
  wire   n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n100, n101;

  DFFR_X1 \Reg_reg[15]  ( .D(n53), .CK(clk), .RN(n54), .Q(dataOut[15]), .QN(
        n70) );
  DFFR_X1 \Reg_reg[14]  ( .D(n55), .CK(clk), .RN(n54), .Q(dataOut[14]), .QN(
        n71) );
  DFFR_X1 \Reg_reg[13]  ( .D(n56), .CK(clk), .RN(n54), .Q(dataOut[13]), .QN(
        n72) );
  DFFR_X1 \Reg_reg[12]  ( .D(n57), .CK(clk), .RN(n54), .Q(dataOut[12]), .QN(
        n73) );
  DFFR_X1 \Reg_reg[11]  ( .D(n58), .CK(clk), .RN(n54), .Q(dataOut[11]), .QN(
        n74) );
  DFFR_X1 \Reg_reg[10]  ( .D(n59), .CK(clk), .RN(n54), .Q(dataOut[10]), .QN(
        n75) );
  DFFR_X1 \Reg_reg[9]  ( .D(n60), .CK(clk), .RN(n54), .Q(dataOut[9]), .QN(n76)
         );
  DFFR_X1 \Reg_reg[8]  ( .D(n61), .CK(clk), .RN(n54), .Q(dataOut[8]), .QN(n77)
         );
  DFFR_X1 \Reg_reg[7]  ( .D(n62), .CK(clk), .RN(n54), .Q(dataOut[7]), .QN(n78)
         );
  DFFR_X1 \Reg_reg[6]  ( .D(n63), .CK(clk), .RN(n54), .Q(dataOut[6]), .QN(n79)
         );
  DFFR_X1 \Reg_reg[5]  ( .D(n64), .CK(clk), .RN(n54), .Q(dataOut[5]), .QN(n80)
         );
  DFFR_X1 \Reg_reg[4]  ( .D(n65), .CK(clk), .RN(n54), .Q(dataOut[4]), .QN(n81)
         );
  DFFR_X1 \Reg_reg[3]  ( .D(n66), .CK(clk), .RN(n54), .Q(dataOut[3]), .QN(n82)
         );
  DFFR_X1 \Reg_reg[2]  ( .D(n67), .CK(clk), .RN(n54), .Q(dataOut[2]), .QN(n83)
         );
  DFFR_X1 \Reg_reg[1]  ( .D(n68), .CK(clk), .RN(n54), .Q(dataOut[1]), .QN(n84)
         );
  DFFR_X1 \Reg_reg[0]  ( .D(n69), .CK(clk), .RN(n54), .Q(dataOut[0]), .QN(n85)
         );
  OAI21_X1 U2 ( .B1(n50), .B2(n85), .A(n101), .ZN(n69) );
  NAND2_X1 U3 ( .A1(n52), .A2(data[0]), .ZN(n101) );
  OAI21_X1 U4 ( .B1(n50), .B2(n84), .A(n100), .ZN(n68) );
  NAND2_X1 U5 ( .A1(data[1]), .A2(n52), .ZN(n100) );
  OAI21_X1 U6 ( .B1(n50), .B2(n83), .A(n99), .ZN(n67) );
  NAND2_X1 U7 ( .A1(data[2]), .A2(n52), .ZN(n99) );
  OAI21_X1 U8 ( .B1(n50), .B2(n82), .A(n98), .ZN(n66) );
  NAND2_X1 U9 ( .A1(data[3]), .A2(n52), .ZN(n98) );
  OAI21_X1 U10 ( .B1(n50), .B2(n81), .A(n97), .ZN(n65) );
  NAND2_X1 U11 ( .A1(data[4]), .A2(n52), .ZN(n97) );
  OAI21_X1 U12 ( .B1(n50), .B2(n80), .A(n96), .ZN(n64) );
  NAND2_X1 U13 ( .A1(data[5]), .A2(n52), .ZN(n96) );
  OAI21_X1 U14 ( .B1(n50), .B2(n79), .A(n95), .ZN(n63) );
  NAND2_X1 U15 ( .A1(data[6]), .A2(n52), .ZN(n95) );
  OAI21_X1 U16 ( .B1(n51), .B2(n78), .A(n94), .ZN(n62) );
  NAND2_X1 U17 ( .A1(data[7]), .A2(n52), .ZN(n94) );
  OAI21_X1 U18 ( .B1(n51), .B2(n77), .A(n93), .ZN(n61) );
  NAND2_X1 U19 ( .A1(data[8]), .A2(n51), .ZN(n93) );
  OAI21_X1 U20 ( .B1(n51), .B2(n76), .A(n92), .ZN(n60) );
  NAND2_X1 U21 ( .A1(data[9]), .A2(n51), .ZN(n92) );
  OAI21_X1 U22 ( .B1(n50), .B2(n75), .A(n91), .ZN(n59) );
  NAND2_X1 U23 ( .A1(data[10]), .A2(n51), .ZN(n91) );
  OAI21_X1 U24 ( .B1(n51), .B2(n74), .A(n90), .ZN(n58) );
  NAND2_X1 U25 ( .A1(data[11]), .A2(n51), .ZN(n90) );
  OAI21_X1 U26 ( .B1(n50), .B2(n73), .A(n89), .ZN(n57) );
  NAND2_X1 U27 ( .A1(data[12]), .A2(n51), .ZN(n89) );
  OAI21_X1 U28 ( .B1(n50), .B2(n72), .A(n88), .ZN(n56) );
  NAND2_X1 U29 ( .A1(data[13]), .A2(n51), .ZN(n88) );
  OAI21_X1 U30 ( .B1(n50), .B2(n71), .A(n87), .ZN(n55) );
  NAND2_X1 U31 ( .A1(data[14]), .A2(n51), .ZN(n87) );
  INV_X1 U32 ( .A(reset), .ZN(n54) );
  OAI21_X1 U33 ( .B1(n50), .B2(n70), .A(n86), .ZN(n53) );
  NAND2_X1 U34 ( .A1(data[15]), .A2(n51), .ZN(n86) );
  CLKBUF_X3 U35 ( .A(write), .Z(n50) );
  CLKBUF_X3 U36 ( .A(write), .Z(n51) );
  CLKBUF_X3 U37 ( .A(write), .Z(n52) );
endmodule


module SingleReg_18 ( data, clk, reset, write, dataOut );
  input [15:0] data;
  output [15:0] dataOut;
  input clk, reset, write;
  wire   n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n100, n101;

  DFFR_X1 \Reg_reg[15]  ( .D(n53), .CK(clk), .RN(n54), .Q(dataOut[15]), .QN(
        n70) );
  DFFR_X1 \Reg_reg[14]  ( .D(n55), .CK(clk), .RN(n54), .Q(dataOut[14]), .QN(
        n71) );
  DFFR_X1 \Reg_reg[13]  ( .D(n56), .CK(clk), .RN(n54), .Q(dataOut[13]), .QN(
        n72) );
  DFFR_X1 \Reg_reg[12]  ( .D(n57), .CK(clk), .RN(n54), .Q(dataOut[12]), .QN(
        n73) );
  DFFR_X1 \Reg_reg[11]  ( .D(n58), .CK(clk), .RN(n54), .Q(dataOut[11]), .QN(
        n74) );
  DFFR_X1 \Reg_reg[10]  ( .D(n59), .CK(clk), .RN(n54), .Q(dataOut[10]), .QN(
        n75) );
  DFFR_X1 \Reg_reg[9]  ( .D(n60), .CK(clk), .RN(n54), .Q(dataOut[9]), .QN(n76)
         );
  DFFR_X1 \Reg_reg[8]  ( .D(n61), .CK(clk), .RN(n54), .Q(dataOut[8]), .QN(n77)
         );
  DFFR_X1 \Reg_reg[7]  ( .D(n62), .CK(clk), .RN(n54), .Q(dataOut[7]), .QN(n78)
         );
  DFFR_X1 \Reg_reg[6]  ( .D(n63), .CK(clk), .RN(n54), .Q(dataOut[6]), .QN(n79)
         );
  DFFR_X1 \Reg_reg[5]  ( .D(n64), .CK(clk), .RN(n54), .Q(dataOut[5]), .QN(n80)
         );
  DFFR_X1 \Reg_reg[4]  ( .D(n65), .CK(clk), .RN(n54), .Q(dataOut[4]), .QN(n81)
         );
  DFFR_X1 \Reg_reg[3]  ( .D(n66), .CK(clk), .RN(n54), .Q(dataOut[3]), .QN(n82)
         );
  DFFR_X1 \Reg_reg[2]  ( .D(n67), .CK(clk), .RN(n54), .Q(dataOut[2]), .QN(n83)
         );
  DFFR_X1 \Reg_reg[1]  ( .D(n68), .CK(clk), .RN(n54), .Q(dataOut[1]), .QN(n84)
         );
  DFFR_X1 \Reg_reg[0]  ( .D(n69), .CK(clk), .RN(n54), .Q(dataOut[0]), .QN(n85)
         );
  OAI21_X1 U2 ( .B1(n50), .B2(n85), .A(n101), .ZN(n69) );
  NAND2_X1 U3 ( .A1(n52), .A2(data[0]), .ZN(n101) );
  OAI21_X1 U4 ( .B1(n50), .B2(n84), .A(n100), .ZN(n68) );
  NAND2_X1 U5 ( .A1(data[1]), .A2(n52), .ZN(n100) );
  OAI21_X1 U6 ( .B1(n50), .B2(n83), .A(n99), .ZN(n67) );
  NAND2_X1 U7 ( .A1(data[2]), .A2(n52), .ZN(n99) );
  OAI21_X1 U8 ( .B1(n50), .B2(n82), .A(n98), .ZN(n66) );
  NAND2_X1 U9 ( .A1(data[3]), .A2(n52), .ZN(n98) );
  OAI21_X1 U10 ( .B1(n50), .B2(n81), .A(n97), .ZN(n65) );
  NAND2_X1 U11 ( .A1(data[4]), .A2(n52), .ZN(n97) );
  OAI21_X1 U12 ( .B1(n50), .B2(n80), .A(n96), .ZN(n64) );
  NAND2_X1 U13 ( .A1(data[5]), .A2(n52), .ZN(n96) );
  OAI21_X1 U14 ( .B1(n50), .B2(n79), .A(n95), .ZN(n63) );
  NAND2_X1 U15 ( .A1(data[6]), .A2(n52), .ZN(n95) );
  OAI21_X1 U16 ( .B1(n51), .B2(n78), .A(n94), .ZN(n62) );
  NAND2_X1 U17 ( .A1(data[7]), .A2(n52), .ZN(n94) );
  OAI21_X1 U18 ( .B1(n51), .B2(n77), .A(n93), .ZN(n61) );
  NAND2_X1 U19 ( .A1(data[8]), .A2(n51), .ZN(n93) );
  OAI21_X1 U20 ( .B1(n51), .B2(n76), .A(n92), .ZN(n60) );
  NAND2_X1 U21 ( .A1(data[9]), .A2(n51), .ZN(n92) );
  OAI21_X1 U22 ( .B1(n50), .B2(n75), .A(n91), .ZN(n59) );
  NAND2_X1 U23 ( .A1(data[10]), .A2(n51), .ZN(n91) );
  OAI21_X1 U24 ( .B1(n51), .B2(n74), .A(n90), .ZN(n58) );
  NAND2_X1 U25 ( .A1(data[11]), .A2(n51), .ZN(n90) );
  OAI21_X1 U26 ( .B1(n50), .B2(n73), .A(n89), .ZN(n57) );
  NAND2_X1 U27 ( .A1(data[12]), .A2(n51), .ZN(n89) );
  OAI21_X1 U28 ( .B1(n50), .B2(n72), .A(n88), .ZN(n56) );
  NAND2_X1 U29 ( .A1(data[13]), .A2(n51), .ZN(n88) );
  OAI21_X1 U30 ( .B1(n50), .B2(n71), .A(n87), .ZN(n55) );
  NAND2_X1 U31 ( .A1(data[14]), .A2(n51), .ZN(n87) );
  INV_X1 U32 ( .A(reset), .ZN(n54) );
  OAI21_X1 U33 ( .B1(n50), .B2(n70), .A(n86), .ZN(n53) );
  NAND2_X1 U34 ( .A1(data[15]), .A2(n51), .ZN(n86) );
  CLKBUF_X3 U35 ( .A(write), .Z(n50) );
  CLKBUF_X3 U36 ( .A(write), .Z(n51) );
  CLKBUF_X3 U37 ( .A(write), .Z(n52) );
endmodule


module SingleReg_17 ( data, clk, reset, write, dataOut );
  input [15:0] data;
  output [15:0] dataOut;
  input clk, reset, write;
  wire   n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n100, n101;

  DFFR_X1 \Reg_reg[15]  ( .D(n53), .CK(clk), .RN(n54), .Q(dataOut[15]), .QN(
        n70) );
  DFFR_X1 \Reg_reg[14]  ( .D(n55), .CK(clk), .RN(n54), .Q(dataOut[14]), .QN(
        n71) );
  DFFR_X1 \Reg_reg[13]  ( .D(n56), .CK(clk), .RN(n54), .Q(dataOut[13]), .QN(
        n72) );
  DFFR_X1 \Reg_reg[12]  ( .D(n57), .CK(clk), .RN(n54), .Q(dataOut[12]), .QN(
        n73) );
  DFFR_X1 \Reg_reg[11]  ( .D(n58), .CK(clk), .RN(n54), .Q(dataOut[11]), .QN(
        n74) );
  DFFR_X1 \Reg_reg[10]  ( .D(n59), .CK(clk), .RN(n54), .Q(dataOut[10]), .QN(
        n75) );
  DFFR_X1 \Reg_reg[9]  ( .D(n60), .CK(clk), .RN(n54), .Q(dataOut[9]), .QN(n76)
         );
  DFFR_X1 \Reg_reg[8]  ( .D(n61), .CK(clk), .RN(n54), .Q(dataOut[8]), .QN(n77)
         );
  DFFR_X1 \Reg_reg[7]  ( .D(n62), .CK(clk), .RN(n54), .Q(dataOut[7]), .QN(n78)
         );
  DFFR_X1 \Reg_reg[6]  ( .D(n63), .CK(clk), .RN(n54), .Q(dataOut[6]), .QN(n79)
         );
  DFFR_X1 \Reg_reg[5]  ( .D(n64), .CK(clk), .RN(n54), .Q(dataOut[5]), .QN(n80)
         );
  DFFR_X1 \Reg_reg[4]  ( .D(n65), .CK(clk), .RN(n54), .Q(dataOut[4]), .QN(n81)
         );
  DFFR_X1 \Reg_reg[3]  ( .D(n66), .CK(clk), .RN(n54), .Q(dataOut[3]), .QN(n82)
         );
  DFFR_X1 \Reg_reg[2]  ( .D(n67), .CK(clk), .RN(n54), .Q(dataOut[2]), .QN(n83)
         );
  DFFR_X1 \Reg_reg[1]  ( .D(n68), .CK(clk), .RN(n54), .Q(dataOut[1]), .QN(n84)
         );
  DFFR_X1 \Reg_reg[0]  ( .D(n69), .CK(clk), .RN(n54), .Q(dataOut[0]), .QN(n85)
         );
  OAI21_X1 U2 ( .B1(n50), .B2(n85), .A(n101), .ZN(n69) );
  NAND2_X1 U3 ( .A1(n52), .A2(data[0]), .ZN(n101) );
  OAI21_X1 U4 ( .B1(n50), .B2(n84), .A(n100), .ZN(n68) );
  NAND2_X1 U5 ( .A1(data[1]), .A2(n52), .ZN(n100) );
  OAI21_X1 U6 ( .B1(n50), .B2(n83), .A(n99), .ZN(n67) );
  NAND2_X1 U7 ( .A1(data[2]), .A2(n52), .ZN(n99) );
  OAI21_X1 U8 ( .B1(n50), .B2(n82), .A(n98), .ZN(n66) );
  NAND2_X1 U9 ( .A1(data[3]), .A2(n52), .ZN(n98) );
  OAI21_X1 U10 ( .B1(n50), .B2(n81), .A(n97), .ZN(n65) );
  NAND2_X1 U11 ( .A1(data[4]), .A2(n52), .ZN(n97) );
  OAI21_X1 U12 ( .B1(n50), .B2(n80), .A(n96), .ZN(n64) );
  NAND2_X1 U13 ( .A1(data[5]), .A2(n52), .ZN(n96) );
  OAI21_X1 U14 ( .B1(n50), .B2(n79), .A(n95), .ZN(n63) );
  NAND2_X1 U15 ( .A1(data[6]), .A2(n52), .ZN(n95) );
  OAI21_X1 U16 ( .B1(n51), .B2(n78), .A(n94), .ZN(n62) );
  NAND2_X1 U17 ( .A1(data[7]), .A2(n52), .ZN(n94) );
  OAI21_X1 U18 ( .B1(n51), .B2(n77), .A(n93), .ZN(n61) );
  NAND2_X1 U19 ( .A1(data[8]), .A2(n51), .ZN(n93) );
  OAI21_X1 U20 ( .B1(n51), .B2(n76), .A(n92), .ZN(n60) );
  NAND2_X1 U21 ( .A1(data[9]), .A2(n51), .ZN(n92) );
  OAI21_X1 U22 ( .B1(n50), .B2(n75), .A(n91), .ZN(n59) );
  NAND2_X1 U23 ( .A1(data[10]), .A2(n51), .ZN(n91) );
  OAI21_X1 U24 ( .B1(n51), .B2(n74), .A(n90), .ZN(n58) );
  NAND2_X1 U25 ( .A1(data[11]), .A2(n51), .ZN(n90) );
  OAI21_X1 U26 ( .B1(n50), .B2(n73), .A(n89), .ZN(n57) );
  NAND2_X1 U27 ( .A1(data[12]), .A2(n51), .ZN(n89) );
  OAI21_X1 U28 ( .B1(n50), .B2(n72), .A(n88), .ZN(n56) );
  NAND2_X1 U29 ( .A1(data[13]), .A2(n51), .ZN(n88) );
  OAI21_X1 U30 ( .B1(n50), .B2(n71), .A(n87), .ZN(n55) );
  NAND2_X1 U31 ( .A1(data[14]), .A2(n51), .ZN(n87) );
  INV_X1 U32 ( .A(reset), .ZN(n54) );
  OAI21_X1 U33 ( .B1(n50), .B2(n70), .A(n86), .ZN(n53) );
  NAND2_X1 U34 ( .A1(data[15]), .A2(n51), .ZN(n86) );
  CLKBUF_X3 U35 ( .A(write), .Z(n50) );
  CLKBUF_X3 U36 ( .A(write), .Z(n51) );
  CLKBUF_X3 U37 ( .A(write), .Z(n52) );
endmodule


module SingleReg_16 ( data, clk, reset, write, dataOut );
  input [15:0] data;
  output [15:0] dataOut;
  input clk, reset, write;
  wire   n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n100, n101;

  DFFR_X1 \Reg_reg[15]  ( .D(n53), .CK(clk), .RN(n54), .Q(dataOut[15]), .QN(
        n70) );
  DFFR_X1 \Reg_reg[14]  ( .D(n55), .CK(clk), .RN(n54), .Q(dataOut[14]), .QN(
        n71) );
  DFFR_X1 \Reg_reg[13]  ( .D(n56), .CK(clk), .RN(n54), .Q(dataOut[13]), .QN(
        n72) );
  DFFR_X1 \Reg_reg[12]  ( .D(n57), .CK(clk), .RN(n54), .Q(dataOut[12]), .QN(
        n73) );
  DFFR_X1 \Reg_reg[11]  ( .D(n58), .CK(clk), .RN(n54), .Q(dataOut[11]), .QN(
        n74) );
  DFFR_X1 \Reg_reg[10]  ( .D(n59), .CK(clk), .RN(n54), .Q(dataOut[10]), .QN(
        n75) );
  DFFR_X1 \Reg_reg[9]  ( .D(n60), .CK(clk), .RN(n54), .Q(dataOut[9]), .QN(n76)
         );
  DFFR_X1 \Reg_reg[8]  ( .D(n61), .CK(clk), .RN(n54), .Q(dataOut[8]), .QN(n77)
         );
  DFFR_X1 \Reg_reg[7]  ( .D(n62), .CK(clk), .RN(n54), .Q(dataOut[7]), .QN(n78)
         );
  DFFR_X1 \Reg_reg[6]  ( .D(n63), .CK(clk), .RN(n54), .Q(dataOut[6]), .QN(n79)
         );
  DFFR_X1 \Reg_reg[5]  ( .D(n64), .CK(clk), .RN(n54), .Q(dataOut[5]), .QN(n80)
         );
  DFFR_X1 \Reg_reg[4]  ( .D(n65), .CK(clk), .RN(n54), .Q(dataOut[4]), .QN(n81)
         );
  DFFR_X1 \Reg_reg[3]  ( .D(n66), .CK(clk), .RN(n54), .Q(dataOut[3]), .QN(n82)
         );
  DFFR_X1 \Reg_reg[2]  ( .D(n67), .CK(clk), .RN(n54), .Q(dataOut[2]), .QN(n83)
         );
  DFFR_X1 \Reg_reg[1]  ( .D(n68), .CK(clk), .RN(n54), .Q(dataOut[1]), .QN(n84)
         );
  DFFR_X1 \Reg_reg[0]  ( .D(n69), .CK(clk), .RN(n54), .Q(dataOut[0]), .QN(n85)
         );
  OAI21_X1 U2 ( .B1(n50), .B2(n85), .A(n101), .ZN(n69) );
  NAND2_X1 U3 ( .A1(n52), .A2(data[0]), .ZN(n101) );
  OAI21_X1 U4 ( .B1(n50), .B2(n84), .A(n100), .ZN(n68) );
  NAND2_X1 U5 ( .A1(data[1]), .A2(n52), .ZN(n100) );
  OAI21_X1 U6 ( .B1(n50), .B2(n83), .A(n99), .ZN(n67) );
  NAND2_X1 U7 ( .A1(data[2]), .A2(n52), .ZN(n99) );
  OAI21_X1 U8 ( .B1(n50), .B2(n82), .A(n98), .ZN(n66) );
  NAND2_X1 U9 ( .A1(data[3]), .A2(n52), .ZN(n98) );
  OAI21_X1 U10 ( .B1(n50), .B2(n81), .A(n97), .ZN(n65) );
  NAND2_X1 U11 ( .A1(data[4]), .A2(n52), .ZN(n97) );
  OAI21_X1 U12 ( .B1(n50), .B2(n80), .A(n96), .ZN(n64) );
  NAND2_X1 U13 ( .A1(data[5]), .A2(n52), .ZN(n96) );
  OAI21_X1 U14 ( .B1(n50), .B2(n79), .A(n95), .ZN(n63) );
  NAND2_X1 U15 ( .A1(data[6]), .A2(n52), .ZN(n95) );
  OAI21_X1 U16 ( .B1(n51), .B2(n78), .A(n94), .ZN(n62) );
  NAND2_X1 U17 ( .A1(data[7]), .A2(n52), .ZN(n94) );
  OAI21_X1 U18 ( .B1(n51), .B2(n77), .A(n93), .ZN(n61) );
  NAND2_X1 U19 ( .A1(data[8]), .A2(n51), .ZN(n93) );
  OAI21_X1 U20 ( .B1(n51), .B2(n76), .A(n92), .ZN(n60) );
  NAND2_X1 U21 ( .A1(data[9]), .A2(n51), .ZN(n92) );
  OAI21_X1 U22 ( .B1(n50), .B2(n75), .A(n91), .ZN(n59) );
  NAND2_X1 U23 ( .A1(data[10]), .A2(n51), .ZN(n91) );
  OAI21_X1 U24 ( .B1(n51), .B2(n74), .A(n90), .ZN(n58) );
  NAND2_X1 U25 ( .A1(data[11]), .A2(n51), .ZN(n90) );
  OAI21_X1 U26 ( .B1(n50), .B2(n73), .A(n89), .ZN(n57) );
  NAND2_X1 U27 ( .A1(data[12]), .A2(n51), .ZN(n89) );
  OAI21_X1 U28 ( .B1(n50), .B2(n72), .A(n88), .ZN(n56) );
  NAND2_X1 U29 ( .A1(data[13]), .A2(n51), .ZN(n88) );
  OAI21_X1 U30 ( .B1(n50), .B2(n71), .A(n87), .ZN(n55) );
  NAND2_X1 U31 ( .A1(data[14]), .A2(n51), .ZN(n87) );
  INV_X1 U32 ( .A(reset), .ZN(n54) );
  OAI21_X1 U33 ( .B1(n50), .B2(n70), .A(n86), .ZN(n53) );
  NAND2_X1 U34 ( .A1(data[15]), .A2(n51), .ZN(n86) );
  CLKBUF_X3 U35 ( .A(write), .Z(n50) );
  CLKBUF_X3 U36 ( .A(write), .Z(n51) );
  CLKBUF_X3 U37 ( .A(write), .Z(n52) );
endmodule


module SingleReg_15 ( data, clk, reset, write, dataOut );
  input [15:0] data;
  output [15:0] dataOut;
  input clk, reset, write;
  wire   n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n100, n101;

  DFFR_X1 \Reg_reg[15]  ( .D(n53), .CK(clk), .RN(n54), .Q(dataOut[15]), .QN(
        n70) );
  DFFR_X1 \Reg_reg[14]  ( .D(n55), .CK(clk), .RN(n54), .Q(dataOut[14]), .QN(
        n71) );
  DFFR_X1 \Reg_reg[13]  ( .D(n56), .CK(clk), .RN(n54), .Q(dataOut[13]), .QN(
        n72) );
  DFFR_X1 \Reg_reg[12]  ( .D(n57), .CK(clk), .RN(n54), .Q(dataOut[12]), .QN(
        n73) );
  DFFR_X1 \Reg_reg[11]  ( .D(n58), .CK(clk), .RN(n54), .Q(dataOut[11]), .QN(
        n74) );
  DFFR_X1 \Reg_reg[10]  ( .D(n59), .CK(clk), .RN(n54), .Q(dataOut[10]), .QN(
        n75) );
  DFFR_X1 \Reg_reg[9]  ( .D(n60), .CK(clk), .RN(n54), .Q(dataOut[9]), .QN(n76)
         );
  DFFR_X1 \Reg_reg[8]  ( .D(n61), .CK(clk), .RN(n54), .Q(dataOut[8]), .QN(n77)
         );
  DFFR_X1 \Reg_reg[7]  ( .D(n62), .CK(clk), .RN(n54), .Q(dataOut[7]), .QN(n78)
         );
  DFFR_X1 \Reg_reg[6]  ( .D(n63), .CK(clk), .RN(n54), .Q(dataOut[6]), .QN(n79)
         );
  DFFR_X1 \Reg_reg[5]  ( .D(n64), .CK(clk), .RN(n54), .Q(dataOut[5]), .QN(n80)
         );
  DFFR_X1 \Reg_reg[4]  ( .D(n65), .CK(clk), .RN(n54), .Q(dataOut[4]), .QN(n81)
         );
  DFFR_X1 \Reg_reg[3]  ( .D(n66), .CK(clk), .RN(n54), .Q(dataOut[3]), .QN(n82)
         );
  DFFR_X1 \Reg_reg[2]  ( .D(n67), .CK(clk), .RN(n54), .Q(dataOut[2]), .QN(n83)
         );
  DFFR_X1 \Reg_reg[1]  ( .D(n68), .CK(clk), .RN(n54), .Q(dataOut[1]), .QN(n84)
         );
  DFFR_X1 \Reg_reg[0]  ( .D(n69), .CK(clk), .RN(n54), .Q(dataOut[0]), .QN(n85)
         );
  OAI21_X1 U2 ( .B1(n50), .B2(n85), .A(n101), .ZN(n69) );
  NAND2_X1 U3 ( .A1(n52), .A2(data[0]), .ZN(n101) );
  OAI21_X1 U4 ( .B1(n50), .B2(n84), .A(n100), .ZN(n68) );
  NAND2_X1 U5 ( .A1(data[1]), .A2(n52), .ZN(n100) );
  OAI21_X1 U6 ( .B1(n50), .B2(n83), .A(n99), .ZN(n67) );
  NAND2_X1 U7 ( .A1(data[2]), .A2(n52), .ZN(n99) );
  OAI21_X1 U8 ( .B1(n50), .B2(n82), .A(n98), .ZN(n66) );
  NAND2_X1 U9 ( .A1(data[3]), .A2(n52), .ZN(n98) );
  OAI21_X1 U10 ( .B1(n50), .B2(n81), .A(n97), .ZN(n65) );
  NAND2_X1 U11 ( .A1(data[4]), .A2(n52), .ZN(n97) );
  OAI21_X1 U12 ( .B1(n50), .B2(n80), .A(n96), .ZN(n64) );
  NAND2_X1 U13 ( .A1(data[5]), .A2(n52), .ZN(n96) );
  OAI21_X1 U14 ( .B1(n50), .B2(n79), .A(n95), .ZN(n63) );
  NAND2_X1 U15 ( .A1(data[6]), .A2(n52), .ZN(n95) );
  OAI21_X1 U16 ( .B1(n51), .B2(n78), .A(n94), .ZN(n62) );
  NAND2_X1 U17 ( .A1(data[7]), .A2(n52), .ZN(n94) );
  OAI21_X1 U18 ( .B1(n51), .B2(n77), .A(n93), .ZN(n61) );
  NAND2_X1 U19 ( .A1(data[8]), .A2(n51), .ZN(n93) );
  OAI21_X1 U20 ( .B1(n51), .B2(n76), .A(n92), .ZN(n60) );
  NAND2_X1 U21 ( .A1(data[9]), .A2(n51), .ZN(n92) );
  OAI21_X1 U22 ( .B1(n50), .B2(n75), .A(n91), .ZN(n59) );
  NAND2_X1 U23 ( .A1(data[10]), .A2(n51), .ZN(n91) );
  OAI21_X1 U24 ( .B1(n51), .B2(n74), .A(n90), .ZN(n58) );
  NAND2_X1 U25 ( .A1(data[11]), .A2(n51), .ZN(n90) );
  OAI21_X1 U26 ( .B1(n50), .B2(n73), .A(n89), .ZN(n57) );
  NAND2_X1 U27 ( .A1(data[12]), .A2(n51), .ZN(n89) );
  OAI21_X1 U28 ( .B1(n50), .B2(n72), .A(n88), .ZN(n56) );
  NAND2_X1 U29 ( .A1(data[13]), .A2(n51), .ZN(n88) );
  OAI21_X1 U30 ( .B1(n50), .B2(n71), .A(n87), .ZN(n55) );
  NAND2_X1 U31 ( .A1(data[14]), .A2(n51), .ZN(n87) );
  INV_X1 U32 ( .A(reset), .ZN(n54) );
  OAI21_X1 U33 ( .B1(n50), .B2(n70), .A(n86), .ZN(n53) );
  NAND2_X1 U34 ( .A1(data[15]), .A2(n51), .ZN(n86) );
  CLKBUF_X3 U35 ( .A(write), .Z(n50) );
  CLKBUF_X3 U36 ( .A(write), .Z(n51) );
  CLKBUF_X3 U37 ( .A(write), .Z(n52) );
endmodule


module SingleReg_14 ( data, clk, reset, write, dataOut );
  input [15:0] data;
  output [15:0] dataOut;
  input clk, reset, write;
  wire   n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n100, n101;

  DFFR_X1 \Reg_reg[15]  ( .D(n53), .CK(clk), .RN(n54), .Q(dataOut[15]), .QN(
        n70) );
  DFFR_X1 \Reg_reg[14]  ( .D(n55), .CK(clk), .RN(n54), .Q(dataOut[14]), .QN(
        n71) );
  DFFR_X1 \Reg_reg[13]  ( .D(n56), .CK(clk), .RN(n54), .Q(dataOut[13]), .QN(
        n72) );
  DFFR_X1 \Reg_reg[12]  ( .D(n57), .CK(clk), .RN(n54), .Q(dataOut[12]), .QN(
        n73) );
  DFFR_X1 \Reg_reg[11]  ( .D(n58), .CK(clk), .RN(n54), .Q(dataOut[11]), .QN(
        n74) );
  DFFR_X1 \Reg_reg[10]  ( .D(n59), .CK(clk), .RN(n54), .Q(dataOut[10]), .QN(
        n75) );
  DFFR_X1 \Reg_reg[9]  ( .D(n60), .CK(clk), .RN(n54), .Q(dataOut[9]), .QN(n76)
         );
  DFFR_X1 \Reg_reg[8]  ( .D(n61), .CK(clk), .RN(n54), .Q(dataOut[8]), .QN(n77)
         );
  DFFR_X1 \Reg_reg[7]  ( .D(n62), .CK(clk), .RN(n54), .Q(dataOut[7]), .QN(n78)
         );
  DFFR_X1 \Reg_reg[6]  ( .D(n63), .CK(clk), .RN(n54), .Q(dataOut[6]), .QN(n79)
         );
  DFFR_X1 \Reg_reg[5]  ( .D(n64), .CK(clk), .RN(n54), .Q(dataOut[5]), .QN(n80)
         );
  DFFR_X1 \Reg_reg[4]  ( .D(n65), .CK(clk), .RN(n54), .Q(dataOut[4]), .QN(n81)
         );
  DFFR_X1 \Reg_reg[3]  ( .D(n66), .CK(clk), .RN(n54), .Q(dataOut[3]), .QN(n82)
         );
  DFFR_X1 \Reg_reg[2]  ( .D(n67), .CK(clk), .RN(n54), .Q(dataOut[2]), .QN(n83)
         );
  DFFR_X1 \Reg_reg[1]  ( .D(n68), .CK(clk), .RN(n54), .Q(dataOut[1]), .QN(n84)
         );
  DFFR_X1 \Reg_reg[0]  ( .D(n69), .CK(clk), .RN(n54), .Q(dataOut[0]), .QN(n85)
         );
  OAI21_X1 U2 ( .B1(n50), .B2(n85), .A(n101), .ZN(n69) );
  NAND2_X1 U3 ( .A1(n52), .A2(data[0]), .ZN(n101) );
  OAI21_X1 U4 ( .B1(n50), .B2(n84), .A(n100), .ZN(n68) );
  NAND2_X1 U5 ( .A1(data[1]), .A2(n52), .ZN(n100) );
  OAI21_X1 U6 ( .B1(n50), .B2(n83), .A(n99), .ZN(n67) );
  NAND2_X1 U7 ( .A1(data[2]), .A2(n52), .ZN(n99) );
  OAI21_X1 U8 ( .B1(n50), .B2(n82), .A(n98), .ZN(n66) );
  NAND2_X1 U9 ( .A1(data[3]), .A2(n52), .ZN(n98) );
  OAI21_X1 U10 ( .B1(n50), .B2(n81), .A(n97), .ZN(n65) );
  NAND2_X1 U11 ( .A1(data[4]), .A2(n52), .ZN(n97) );
  OAI21_X1 U12 ( .B1(n50), .B2(n80), .A(n96), .ZN(n64) );
  NAND2_X1 U13 ( .A1(data[5]), .A2(n52), .ZN(n96) );
  OAI21_X1 U14 ( .B1(n50), .B2(n79), .A(n95), .ZN(n63) );
  NAND2_X1 U15 ( .A1(data[6]), .A2(n52), .ZN(n95) );
  OAI21_X1 U16 ( .B1(n51), .B2(n78), .A(n94), .ZN(n62) );
  NAND2_X1 U17 ( .A1(data[7]), .A2(n52), .ZN(n94) );
  OAI21_X1 U18 ( .B1(n51), .B2(n77), .A(n93), .ZN(n61) );
  NAND2_X1 U19 ( .A1(data[8]), .A2(n51), .ZN(n93) );
  OAI21_X1 U20 ( .B1(n51), .B2(n76), .A(n92), .ZN(n60) );
  NAND2_X1 U21 ( .A1(data[9]), .A2(n51), .ZN(n92) );
  OAI21_X1 U22 ( .B1(n50), .B2(n75), .A(n91), .ZN(n59) );
  NAND2_X1 U23 ( .A1(data[10]), .A2(n51), .ZN(n91) );
  OAI21_X1 U24 ( .B1(n51), .B2(n74), .A(n90), .ZN(n58) );
  NAND2_X1 U25 ( .A1(data[11]), .A2(n51), .ZN(n90) );
  OAI21_X1 U26 ( .B1(n50), .B2(n73), .A(n89), .ZN(n57) );
  NAND2_X1 U27 ( .A1(data[12]), .A2(n51), .ZN(n89) );
  OAI21_X1 U28 ( .B1(n50), .B2(n72), .A(n88), .ZN(n56) );
  NAND2_X1 U29 ( .A1(data[13]), .A2(n51), .ZN(n88) );
  OAI21_X1 U30 ( .B1(n50), .B2(n71), .A(n87), .ZN(n55) );
  NAND2_X1 U31 ( .A1(data[14]), .A2(n51), .ZN(n87) );
  INV_X1 U32 ( .A(reset), .ZN(n54) );
  OAI21_X1 U33 ( .B1(n50), .B2(n70), .A(n86), .ZN(n53) );
  NAND2_X1 U34 ( .A1(data[15]), .A2(n51), .ZN(n86) );
  CLKBUF_X3 U35 ( .A(write), .Z(n50) );
  CLKBUF_X3 U36 ( .A(write), .Z(n51) );
  CLKBUF_X3 U37 ( .A(write), .Z(n52) );
endmodule


module SingleReg_13 ( data, clk, reset, write, dataOut );
  input [15:0] data;
  output [15:0] dataOut;
  input clk, reset, write;
  wire   n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n100, n101;

  DFFR_X1 \Reg_reg[15]  ( .D(n53), .CK(clk), .RN(n54), .Q(dataOut[15]), .QN(
        n70) );
  DFFR_X1 \Reg_reg[14]  ( .D(n55), .CK(clk), .RN(n54), .Q(dataOut[14]), .QN(
        n71) );
  DFFR_X1 \Reg_reg[13]  ( .D(n56), .CK(clk), .RN(n54), .Q(dataOut[13]), .QN(
        n72) );
  DFFR_X1 \Reg_reg[12]  ( .D(n57), .CK(clk), .RN(n54), .Q(dataOut[12]), .QN(
        n73) );
  DFFR_X1 \Reg_reg[11]  ( .D(n58), .CK(clk), .RN(n54), .Q(dataOut[11]), .QN(
        n74) );
  DFFR_X1 \Reg_reg[10]  ( .D(n59), .CK(clk), .RN(n54), .Q(dataOut[10]), .QN(
        n75) );
  DFFR_X1 \Reg_reg[9]  ( .D(n60), .CK(clk), .RN(n54), .Q(dataOut[9]), .QN(n76)
         );
  DFFR_X1 \Reg_reg[8]  ( .D(n61), .CK(clk), .RN(n54), .Q(dataOut[8]), .QN(n77)
         );
  DFFR_X1 \Reg_reg[7]  ( .D(n62), .CK(clk), .RN(n54), .Q(dataOut[7]), .QN(n78)
         );
  DFFR_X1 \Reg_reg[6]  ( .D(n63), .CK(clk), .RN(n54), .Q(dataOut[6]), .QN(n79)
         );
  DFFR_X1 \Reg_reg[5]  ( .D(n64), .CK(clk), .RN(n54), .Q(dataOut[5]), .QN(n80)
         );
  DFFR_X1 \Reg_reg[4]  ( .D(n65), .CK(clk), .RN(n54), .Q(dataOut[4]), .QN(n81)
         );
  DFFR_X1 \Reg_reg[3]  ( .D(n66), .CK(clk), .RN(n54), .Q(dataOut[3]), .QN(n82)
         );
  DFFR_X1 \Reg_reg[2]  ( .D(n67), .CK(clk), .RN(n54), .Q(dataOut[2]), .QN(n83)
         );
  DFFR_X1 \Reg_reg[1]  ( .D(n68), .CK(clk), .RN(n54), .Q(dataOut[1]), .QN(n84)
         );
  DFFR_X1 \Reg_reg[0]  ( .D(n69), .CK(clk), .RN(n54), .Q(dataOut[0]), .QN(n85)
         );
  OAI21_X1 U2 ( .B1(n50), .B2(n85), .A(n101), .ZN(n69) );
  NAND2_X1 U3 ( .A1(n52), .A2(data[0]), .ZN(n101) );
  OAI21_X1 U4 ( .B1(n50), .B2(n84), .A(n100), .ZN(n68) );
  NAND2_X1 U5 ( .A1(data[1]), .A2(n52), .ZN(n100) );
  OAI21_X1 U6 ( .B1(n50), .B2(n83), .A(n99), .ZN(n67) );
  NAND2_X1 U7 ( .A1(data[2]), .A2(n52), .ZN(n99) );
  OAI21_X1 U8 ( .B1(n50), .B2(n82), .A(n98), .ZN(n66) );
  NAND2_X1 U9 ( .A1(data[3]), .A2(n52), .ZN(n98) );
  OAI21_X1 U10 ( .B1(n50), .B2(n81), .A(n97), .ZN(n65) );
  NAND2_X1 U11 ( .A1(data[4]), .A2(n52), .ZN(n97) );
  OAI21_X1 U12 ( .B1(n50), .B2(n80), .A(n96), .ZN(n64) );
  NAND2_X1 U13 ( .A1(data[5]), .A2(n52), .ZN(n96) );
  OAI21_X1 U14 ( .B1(n50), .B2(n79), .A(n95), .ZN(n63) );
  NAND2_X1 U15 ( .A1(data[6]), .A2(n52), .ZN(n95) );
  OAI21_X1 U16 ( .B1(n51), .B2(n78), .A(n94), .ZN(n62) );
  NAND2_X1 U17 ( .A1(data[7]), .A2(n52), .ZN(n94) );
  OAI21_X1 U18 ( .B1(n51), .B2(n77), .A(n93), .ZN(n61) );
  NAND2_X1 U19 ( .A1(data[8]), .A2(n51), .ZN(n93) );
  OAI21_X1 U20 ( .B1(n51), .B2(n76), .A(n92), .ZN(n60) );
  NAND2_X1 U21 ( .A1(data[9]), .A2(n51), .ZN(n92) );
  OAI21_X1 U22 ( .B1(n50), .B2(n75), .A(n91), .ZN(n59) );
  NAND2_X1 U23 ( .A1(data[10]), .A2(n51), .ZN(n91) );
  OAI21_X1 U24 ( .B1(n51), .B2(n74), .A(n90), .ZN(n58) );
  NAND2_X1 U25 ( .A1(data[11]), .A2(n51), .ZN(n90) );
  OAI21_X1 U26 ( .B1(n50), .B2(n73), .A(n89), .ZN(n57) );
  NAND2_X1 U27 ( .A1(data[12]), .A2(n51), .ZN(n89) );
  OAI21_X1 U28 ( .B1(n50), .B2(n72), .A(n88), .ZN(n56) );
  NAND2_X1 U29 ( .A1(data[13]), .A2(n51), .ZN(n88) );
  OAI21_X1 U30 ( .B1(n50), .B2(n71), .A(n87), .ZN(n55) );
  NAND2_X1 U31 ( .A1(data[14]), .A2(n51), .ZN(n87) );
  INV_X1 U32 ( .A(reset), .ZN(n54) );
  OAI21_X1 U33 ( .B1(n50), .B2(n70), .A(n86), .ZN(n53) );
  NAND2_X1 U34 ( .A1(data[15]), .A2(n51), .ZN(n86) );
  CLKBUF_X3 U35 ( .A(write), .Z(n50) );
  CLKBUF_X3 U36 ( .A(write), .Z(n51) );
  CLKBUF_X3 U37 ( .A(write), .Z(n52) );
endmodule


module SingleReg_12 ( data, clk, reset, write, dataOut );
  input [15:0] data;
  output [15:0] dataOut;
  input clk, reset, write;
  wire   n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n100, n101;

  DFFR_X1 \Reg_reg[15]  ( .D(n53), .CK(clk), .RN(n54), .Q(dataOut[15]), .QN(
        n70) );
  DFFR_X1 \Reg_reg[14]  ( .D(n55), .CK(clk), .RN(n54), .Q(dataOut[14]), .QN(
        n71) );
  DFFR_X1 \Reg_reg[13]  ( .D(n56), .CK(clk), .RN(n54), .Q(dataOut[13]), .QN(
        n72) );
  DFFR_X1 \Reg_reg[12]  ( .D(n57), .CK(clk), .RN(n54), .Q(dataOut[12]), .QN(
        n73) );
  DFFR_X1 \Reg_reg[11]  ( .D(n58), .CK(clk), .RN(n54), .Q(dataOut[11]), .QN(
        n74) );
  DFFR_X1 \Reg_reg[10]  ( .D(n59), .CK(clk), .RN(n54), .Q(dataOut[10]), .QN(
        n75) );
  DFFR_X1 \Reg_reg[9]  ( .D(n60), .CK(clk), .RN(n54), .Q(dataOut[9]), .QN(n76)
         );
  DFFR_X1 \Reg_reg[8]  ( .D(n61), .CK(clk), .RN(n54), .Q(dataOut[8]), .QN(n77)
         );
  DFFR_X1 \Reg_reg[7]  ( .D(n62), .CK(clk), .RN(n54), .Q(dataOut[7]), .QN(n78)
         );
  DFFR_X1 \Reg_reg[6]  ( .D(n63), .CK(clk), .RN(n54), .Q(dataOut[6]), .QN(n79)
         );
  DFFR_X1 \Reg_reg[5]  ( .D(n64), .CK(clk), .RN(n54), .Q(dataOut[5]), .QN(n80)
         );
  DFFR_X1 \Reg_reg[4]  ( .D(n65), .CK(clk), .RN(n54), .Q(dataOut[4]), .QN(n81)
         );
  DFFR_X1 \Reg_reg[3]  ( .D(n66), .CK(clk), .RN(n54), .Q(dataOut[3]), .QN(n82)
         );
  DFFR_X1 \Reg_reg[2]  ( .D(n67), .CK(clk), .RN(n54), .Q(dataOut[2]), .QN(n83)
         );
  DFFR_X1 \Reg_reg[1]  ( .D(n68), .CK(clk), .RN(n54), .Q(dataOut[1]), .QN(n84)
         );
  DFFR_X1 \Reg_reg[0]  ( .D(n69), .CK(clk), .RN(n54), .Q(dataOut[0]), .QN(n85)
         );
  OAI21_X1 U2 ( .B1(n50), .B2(n85), .A(n101), .ZN(n69) );
  NAND2_X1 U3 ( .A1(n52), .A2(data[0]), .ZN(n101) );
  OAI21_X1 U4 ( .B1(n50), .B2(n84), .A(n100), .ZN(n68) );
  NAND2_X1 U5 ( .A1(data[1]), .A2(n52), .ZN(n100) );
  OAI21_X1 U6 ( .B1(n50), .B2(n83), .A(n99), .ZN(n67) );
  NAND2_X1 U7 ( .A1(data[2]), .A2(n52), .ZN(n99) );
  OAI21_X1 U8 ( .B1(n50), .B2(n82), .A(n98), .ZN(n66) );
  NAND2_X1 U9 ( .A1(data[3]), .A2(n52), .ZN(n98) );
  OAI21_X1 U10 ( .B1(n50), .B2(n81), .A(n97), .ZN(n65) );
  NAND2_X1 U11 ( .A1(data[4]), .A2(n52), .ZN(n97) );
  OAI21_X1 U12 ( .B1(n50), .B2(n80), .A(n96), .ZN(n64) );
  NAND2_X1 U13 ( .A1(data[5]), .A2(n52), .ZN(n96) );
  OAI21_X1 U14 ( .B1(n50), .B2(n79), .A(n95), .ZN(n63) );
  NAND2_X1 U15 ( .A1(data[6]), .A2(n52), .ZN(n95) );
  OAI21_X1 U16 ( .B1(n51), .B2(n78), .A(n94), .ZN(n62) );
  NAND2_X1 U17 ( .A1(data[7]), .A2(n52), .ZN(n94) );
  OAI21_X1 U18 ( .B1(n51), .B2(n77), .A(n93), .ZN(n61) );
  NAND2_X1 U19 ( .A1(data[8]), .A2(n51), .ZN(n93) );
  OAI21_X1 U20 ( .B1(n51), .B2(n76), .A(n92), .ZN(n60) );
  NAND2_X1 U21 ( .A1(data[9]), .A2(n51), .ZN(n92) );
  OAI21_X1 U22 ( .B1(n50), .B2(n75), .A(n91), .ZN(n59) );
  NAND2_X1 U23 ( .A1(data[10]), .A2(n51), .ZN(n91) );
  OAI21_X1 U24 ( .B1(n51), .B2(n74), .A(n90), .ZN(n58) );
  NAND2_X1 U25 ( .A1(data[11]), .A2(n51), .ZN(n90) );
  OAI21_X1 U26 ( .B1(n50), .B2(n73), .A(n89), .ZN(n57) );
  NAND2_X1 U27 ( .A1(data[12]), .A2(n51), .ZN(n89) );
  OAI21_X1 U28 ( .B1(n50), .B2(n72), .A(n88), .ZN(n56) );
  NAND2_X1 U29 ( .A1(data[13]), .A2(n51), .ZN(n88) );
  OAI21_X1 U30 ( .B1(n50), .B2(n71), .A(n87), .ZN(n55) );
  NAND2_X1 U31 ( .A1(data[14]), .A2(n51), .ZN(n87) );
  INV_X1 U32 ( .A(reset), .ZN(n54) );
  OAI21_X1 U33 ( .B1(n50), .B2(n70), .A(n86), .ZN(n53) );
  NAND2_X1 U34 ( .A1(data[15]), .A2(n51), .ZN(n86) );
  CLKBUF_X3 U35 ( .A(write), .Z(n50) );
  CLKBUF_X3 U36 ( .A(write), .Z(n51) );
  CLKBUF_X3 U37 ( .A(write), .Z(n52) );
endmodule


module SingleReg_11 ( data, clk, reset, write, dataOut );
  input [15:0] data;
  output [15:0] dataOut;
  input clk, reset, write;
  wire   n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n100, n101;

  DFFR_X1 \Reg_reg[15]  ( .D(n53), .CK(clk), .RN(n54), .Q(dataOut[15]), .QN(
        n70) );
  DFFR_X1 \Reg_reg[14]  ( .D(n55), .CK(clk), .RN(n54), .Q(dataOut[14]), .QN(
        n71) );
  DFFR_X1 \Reg_reg[13]  ( .D(n56), .CK(clk), .RN(n54), .Q(dataOut[13]), .QN(
        n72) );
  DFFR_X1 \Reg_reg[12]  ( .D(n57), .CK(clk), .RN(n54), .Q(dataOut[12]), .QN(
        n73) );
  DFFR_X1 \Reg_reg[11]  ( .D(n58), .CK(clk), .RN(n54), .Q(dataOut[11]), .QN(
        n74) );
  DFFR_X1 \Reg_reg[10]  ( .D(n59), .CK(clk), .RN(n54), .Q(dataOut[10]), .QN(
        n75) );
  DFFR_X1 \Reg_reg[9]  ( .D(n60), .CK(clk), .RN(n54), .Q(dataOut[9]), .QN(n76)
         );
  DFFR_X1 \Reg_reg[8]  ( .D(n61), .CK(clk), .RN(n54), .Q(dataOut[8]), .QN(n77)
         );
  DFFR_X1 \Reg_reg[7]  ( .D(n62), .CK(clk), .RN(n54), .Q(dataOut[7]), .QN(n78)
         );
  DFFR_X1 \Reg_reg[6]  ( .D(n63), .CK(clk), .RN(n54), .Q(dataOut[6]), .QN(n79)
         );
  DFFR_X1 \Reg_reg[5]  ( .D(n64), .CK(clk), .RN(n54), .Q(dataOut[5]), .QN(n80)
         );
  DFFR_X1 \Reg_reg[4]  ( .D(n65), .CK(clk), .RN(n54), .Q(dataOut[4]), .QN(n81)
         );
  DFFR_X1 \Reg_reg[3]  ( .D(n66), .CK(clk), .RN(n54), .Q(dataOut[3]), .QN(n82)
         );
  DFFR_X1 \Reg_reg[2]  ( .D(n67), .CK(clk), .RN(n54), .Q(dataOut[2]), .QN(n83)
         );
  DFFR_X1 \Reg_reg[1]  ( .D(n68), .CK(clk), .RN(n54), .Q(dataOut[1]), .QN(n84)
         );
  DFFR_X1 \Reg_reg[0]  ( .D(n69), .CK(clk), .RN(n54), .Q(dataOut[0]), .QN(n85)
         );
  OAI21_X1 U2 ( .B1(n50), .B2(n85), .A(n101), .ZN(n69) );
  NAND2_X1 U3 ( .A1(n52), .A2(data[0]), .ZN(n101) );
  OAI21_X1 U4 ( .B1(n50), .B2(n84), .A(n100), .ZN(n68) );
  NAND2_X1 U5 ( .A1(data[1]), .A2(n52), .ZN(n100) );
  OAI21_X1 U6 ( .B1(n50), .B2(n83), .A(n99), .ZN(n67) );
  NAND2_X1 U7 ( .A1(data[2]), .A2(n52), .ZN(n99) );
  OAI21_X1 U8 ( .B1(n50), .B2(n82), .A(n98), .ZN(n66) );
  NAND2_X1 U9 ( .A1(data[3]), .A2(n52), .ZN(n98) );
  OAI21_X1 U10 ( .B1(n50), .B2(n81), .A(n97), .ZN(n65) );
  NAND2_X1 U11 ( .A1(data[4]), .A2(n52), .ZN(n97) );
  OAI21_X1 U12 ( .B1(n50), .B2(n80), .A(n96), .ZN(n64) );
  NAND2_X1 U13 ( .A1(data[5]), .A2(n52), .ZN(n96) );
  OAI21_X1 U14 ( .B1(n50), .B2(n79), .A(n95), .ZN(n63) );
  NAND2_X1 U15 ( .A1(data[6]), .A2(n52), .ZN(n95) );
  OAI21_X1 U16 ( .B1(n51), .B2(n78), .A(n94), .ZN(n62) );
  NAND2_X1 U17 ( .A1(data[7]), .A2(n52), .ZN(n94) );
  OAI21_X1 U18 ( .B1(n51), .B2(n77), .A(n93), .ZN(n61) );
  NAND2_X1 U19 ( .A1(data[8]), .A2(n51), .ZN(n93) );
  OAI21_X1 U20 ( .B1(n51), .B2(n76), .A(n92), .ZN(n60) );
  NAND2_X1 U21 ( .A1(data[9]), .A2(n51), .ZN(n92) );
  OAI21_X1 U22 ( .B1(n50), .B2(n75), .A(n91), .ZN(n59) );
  NAND2_X1 U23 ( .A1(data[10]), .A2(n51), .ZN(n91) );
  OAI21_X1 U24 ( .B1(n51), .B2(n74), .A(n90), .ZN(n58) );
  NAND2_X1 U25 ( .A1(data[11]), .A2(n51), .ZN(n90) );
  OAI21_X1 U26 ( .B1(n50), .B2(n73), .A(n89), .ZN(n57) );
  NAND2_X1 U27 ( .A1(data[12]), .A2(n51), .ZN(n89) );
  OAI21_X1 U28 ( .B1(n50), .B2(n72), .A(n88), .ZN(n56) );
  NAND2_X1 U29 ( .A1(data[13]), .A2(n51), .ZN(n88) );
  OAI21_X1 U30 ( .B1(n50), .B2(n71), .A(n87), .ZN(n55) );
  NAND2_X1 U31 ( .A1(data[14]), .A2(n51), .ZN(n87) );
  INV_X1 U32 ( .A(reset), .ZN(n54) );
  OAI21_X1 U33 ( .B1(n50), .B2(n70), .A(n86), .ZN(n53) );
  NAND2_X1 U34 ( .A1(data[15]), .A2(n51), .ZN(n86) );
  CLKBUF_X3 U35 ( .A(write), .Z(n50) );
  CLKBUF_X3 U36 ( .A(write), .Z(n51) );
  CLKBUF_X3 U37 ( .A(write), .Z(n52) );
endmodule


module SingleReg_10 ( data, clk, reset, write, dataOut );
  input [15:0] data;
  output [15:0] dataOut;
  input clk, reset, write;
  wire   n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n100, n101;

  DFFR_X1 \Reg_reg[15]  ( .D(n53), .CK(clk), .RN(n54), .Q(dataOut[15]), .QN(
        n70) );
  DFFR_X1 \Reg_reg[14]  ( .D(n55), .CK(clk), .RN(n54), .Q(dataOut[14]), .QN(
        n71) );
  DFFR_X1 \Reg_reg[13]  ( .D(n56), .CK(clk), .RN(n54), .Q(dataOut[13]), .QN(
        n72) );
  DFFR_X1 \Reg_reg[12]  ( .D(n57), .CK(clk), .RN(n54), .Q(dataOut[12]), .QN(
        n73) );
  DFFR_X1 \Reg_reg[11]  ( .D(n58), .CK(clk), .RN(n54), .Q(dataOut[11]), .QN(
        n74) );
  DFFR_X1 \Reg_reg[10]  ( .D(n59), .CK(clk), .RN(n54), .Q(dataOut[10]), .QN(
        n75) );
  DFFR_X1 \Reg_reg[9]  ( .D(n60), .CK(clk), .RN(n54), .Q(dataOut[9]), .QN(n76)
         );
  DFFR_X1 \Reg_reg[8]  ( .D(n61), .CK(clk), .RN(n54), .Q(dataOut[8]), .QN(n77)
         );
  DFFR_X1 \Reg_reg[7]  ( .D(n62), .CK(clk), .RN(n54), .Q(dataOut[7]), .QN(n78)
         );
  DFFR_X1 \Reg_reg[6]  ( .D(n63), .CK(clk), .RN(n54), .Q(dataOut[6]), .QN(n79)
         );
  DFFR_X1 \Reg_reg[5]  ( .D(n64), .CK(clk), .RN(n54), .Q(dataOut[5]), .QN(n80)
         );
  DFFR_X1 \Reg_reg[4]  ( .D(n65), .CK(clk), .RN(n54), .Q(dataOut[4]), .QN(n81)
         );
  DFFR_X1 \Reg_reg[3]  ( .D(n66), .CK(clk), .RN(n54), .Q(dataOut[3]), .QN(n82)
         );
  DFFR_X1 \Reg_reg[2]  ( .D(n67), .CK(clk), .RN(n54), .Q(dataOut[2]), .QN(n83)
         );
  DFFR_X1 \Reg_reg[1]  ( .D(n68), .CK(clk), .RN(n54), .Q(dataOut[1]), .QN(n84)
         );
  DFFR_X1 \Reg_reg[0]  ( .D(n69), .CK(clk), .RN(n54), .Q(dataOut[0]), .QN(n85)
         );
  OAI21_X1 U2 ( .B1(n50), .B2(n85), .A(n101), .ZN(n69) );
  NAND2_X1 U3 ( .A1(n52), .A2(data[0]), .ZN(n101) );
  OAI21_X1 U4 ( .B1(n50), .B2(n84), .A(n100), .ZN(n68) );
  NAND2_X1 U5 ( .A1(data[1]), .A2(n52), .ZN(n100) );
  OAI21_X1 U6 ( .B1(n50), .B2(n83), .A(n99), .ZN(n67) );
  NAND2_X1 U7 ( .A1(data[2]), .A2(n52), .ZN(n99) );
  OAI21_X1 U8 ( .B1(n50), .B2(n82), .A(n98), .ZN(n66) );
  NAND2_X1 U9 ( .A1(data[3]), .A2(n52), .ZN(n98) );
  OAI21_X1 U10 ( .B1(n50), .B2(n81), .A(n97), .ZN(n65) );
  NAND2_X1 U11 ( .A1(data[4]), .A2(n52), .ZN(n97) );
  OAI21_X1 U12 ( .B1(n50), .B2(n80), .A(n96), .ZN(n64) );
  NAND2_X1 U13 ( .A1(data[5]), .A2(n52), .ZN(n96) );
  OAI21_X1 U14 ( .B1(n50), .B2(n79), .A(n95), .ZN(n63) );
  NAND2_X1 U15 ( .A1(data[6]), .A2(n52), .ZN(n95) );
  OAI21_X1 U16 ( .B1(n51), .B2(n78), .A(n94), .ZN(n62) );
  NAND2_X1 U17 ( .A1(data[7]), .A2(n52), .ZN(n94) );
  OAI21_X1 U18 ( .B1(n51), .B2(n77), .A(n93), .ZN(n61) );
  NAND2_X1 U19 ( .A1(data[8]), .A2(n51), .ZN(n93) );
  OAI21_X1 U20 ( .B1(n51), .B2(n76), .A(n92), .ZN(n60) );
  NAND2_X1 U21 ( .A1(data[9]), .A2(n51), .ZN(n92) );
  OAI21_X1 U22 ( .B1(n50), .B2(n75), .A(n91), .ZN(n59) );
  NAND2_X1 U23 ( .A1(data[10]), .A2(n51), .ZN(n91) );
  OAI21_X1 U24 ( .B1(n51), .B2(n74), .A(n90), .ZN(n58) );
  NAND2_X1 U25 ( .A1(data[11]), .A2(n51), .ZN(n90) );
  OAI21_X1 U26 ( .B1(n50), .B2(n73), .A(n89), .ZN(n57) );
  NAND2_X1 U27 ( .A1(data[12]), .A2(n51), .ZN(n89) );
  OAI21_X1 U28 ( .B1(n50), .B2(n72), .A(n88), .ZN(n56) );
  NAND2_X1 U29 ( .A1(data[13]), .A2(n51), .ZN(n88) );
  OAI21_X1 U30 ( .B1(n50), .B2(n71), .A(n87), .ZN(n55) );
  NAND2_X1 U31 ( .A1(data[14]), .A2(n51), .ZN(n87) );
  INV_X1 U32 ( .A(reset), .ZN(n54) );
  OAI21_X1 U33 ( .B1(n50), .B2(n70), .A(n86), .ZN(n53) );
  NAND2_X1 U34 ( .A1(data[15]), .A2(n51), .ZN(n86) );
  CLKBUF_X3 U35 ( .A(write), .Z(n50) );
  CLKBUF_X3 U36 ( .A(write), .Z(n51) );
  CLKBUF_X3 U37 ( .A(write), .Z(n52) );
endmodule


module SingleReg_9 ( data, clk, reset, write, dataOut );
  input [15:0] data;
  output [15:0] dataOut;
  input clk, reset, write;
  wire   n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n100, n101;

  DFFR_X1 \Reg_reg[15]  ( .D(n53), .CK(clk), .RN(n54), .Q(dataOut[15]), .QN(
        n70) );
  DFFR_X1 \Reg_reg[14]  ( .D(n55), .CK(clk), .RN(n54), .Q(dataOut[14]), .QN(
        n71) );
  DFFR_X1 \Reg_reg[13]  ( .D(n56), .CK(clk), .RN(n54), .Q(dataOut[13]), .QN(
        n72) );
  DFFR_X1 \Reg_reg[12]  ( .D(n57), .CK(clk), .RN(n54), .Q(dataOut[12]), .QN(
        n73) );
  DFFR_X1 \Reg_reg[11]  ( .D(n58), .CK(clk), .RN(n54), .Q(dataOut[11]), .QN(
        n74) );
  DFFR_X1 \Reg_reg[10]  ( .D(n59), .CK(clk), .RN(n54), .Q(dataOut[10]), .QN(
        n75) );
  DFFR_X1 \Reg_reg[9]  ( .D(n60), .CK(clk), .RN(n54), .Q(dataOut[9]), .QN(n76)
         );
  DFFR_X1 \Reg_reg[8]  ( .D(n61), .CK(clk), .RN(n54), .Q(dataOut[8]), .QN(n77)
         );
  DFFR_X1 \Reg_reg[7]  ( .D(n62), .CK(clk), .RN(n54), .Q(dataOut[7]), .QN(n78)
         );
  DFFR_X1 \Reg_reg[6]  ( .D(n63), .CK(clk), .RN(n54), .Q(dataOut[6]), .QN(n79)
         );
  DFFR_X1 \Reg_reg[5]  ( .D(n64), .CK(clk), .RN(n54), .Q(dataOut[5]), .QN(n80)
         );
  DFFR_X1 \Reg_reg[4]  ( .D(n65), .CK(clk), .RN(n54), .Q(dataOut[4]), .QN(n81)
         );
  DFFR_X1 \Reg_reg[3]  ( .D(n66), .CK(clk), .RN(n54), .Q(dataOut[3]), .QN(n82)
         );
  DFFR_X1 \Reg_reg[2]  ( .D(n67), .CK(clk), .RN(n54), .Q(dataOut[2]), .QN(n83)
         );
  DFFR_X1 \Reg_reg[1]  ( .D(n68), .CK(clk), .RN(n54), .Q(dataOut[1]), .QN(n84)
         );
  DFFR_X1 \Reg_reg[0]  ( .D(n69), .CK(clk), .RN(n54), .Q(dataOut[0]), .QN(n85)
         );
  OAI21_X1 U2 ( .B1(n50), .B2(n85), .A(n101), .ZN(n69) );
  NAND2_X1 U3 ( .A1(n52), .A2(data[0]), .ZN(n101) );
  OAI21_X1 U4 ( .B1(n50), .B2(n84), .A(n100), .ZN(n68) );
  NAND2_X1 U5 ( .A1(data[1]), .A2(n52), .ZN(n100) );
  OAI21_X1 U6 ( .B1(n50), .B2(n83), .A(n99), .ZN(n67) );
  NAND2_X1 U7 ( .A1(data[2]), .A2(n52), .ZN(n99) );
  OAI21_X1 U8 ( .B1(n50), .B2(n82), .A(n98), .ZN(n66) );
  NAND2_X1 U9 ( .A1(data[3]), .A2(n52), .ZN(n98) );
  OAI21_X1 U10 ( .B1(n50), .B2(n81), .A(n97), .ZN(n65) );
  NAND2_X1 U11 ( .A1(data[4]), .A2(n52), .ZN(n97) );
  OAI21_X1 U12 ( .B1(n50), .B2(n80), .A(n96), .ZN(n64) );
  NAND2_X1 U13 ( .A1(data[5]), .A2(n52), .ZN(n96) );
  OAI21_X1 U14 ( .B1(n50), .B2(n79), .A(n95), .ZN(n63) );
  NAND2_X1 U15 ( .A1(data[6]), .A2(n52), .ZN(n95) );
  OAI21_X1 U16 ( .B1(n51), .B2(n78), .A(n94), .ZN(n62) );
  NAND2_X1 U17 ( .A1(data[7]), .A2(n52), .ZN(n94) );
  OAI21_X1 U18 ( .B1(n51), .B2(n77), .A(n93), .ZN(n61) );
  NAND2_X1 U19 ( .A1(data[8]), .A2(n51), .ZN(n93) );
  OAI21_X1 U20 ( .B1(n51), .B2(n76), .A(n92), .ZN(n60) );
  NAND2_X1 U21 ( .A1(data[9]), .A2(n51), .ZN(n92) );
  OAI21_X1 U22 ( .B1(n50), .B2(n75), .A(n91), .ZN(n59) );
  NAND2_X1 U23 ( .A1(data[10]), .A2(n51), .ZN(n91) );
  OAI21_X1 U24 ( .B1(n51), .B2(n74), .A(n90), .ZN(n58) );
  NAND2_X1 U25 ( .A1(data[11]), .A2(n51), .ZN(n90) );
  OAI21_X1 U26 ( .B1(n50), .B2(n73), .A(n89), .ZN(n57) );
  NAND2_X1 U27 ( .A1(data[12]), .A2(n51), .ZN(n89) );
  OAI21_X1 U28 ( .B1(n50), .B2(n72), .A(n88), .ZN(n56) );
  NAND2_X1 U29 ( .A1(data[13]), .A2(n51), .ZN(n88) );
  OAI21_X1 U30 ( .B1(n50), .B2(n71), .A(n87), .ZN(n55) );
  NAND2_X1 U31 ( .A1(data[14]), .A2(n51), .ZN(n87) );
  INV_X1 U32 ( .A(reset), .ZN(n54) );
  OAI21_X1 U33 ( .B1(n50), .B2(n70), .A(n86), .ZN(n53) );
  NAND2_X1 U34 ( .A1(data[15]), .A2(n51), .ZN(n86) );
  CLKBUF_X3 U35 ( .A(write), .Z(n50) );
  CLKBUF_X3 U36 ( .A(write), .Z(n51) );
  CLKBUF_X3 U37 ( .A(write), .Z(n52) );
endmodule


module SingleReg_8 ( data, clk, reset, write, dataOut );
  input [15:0] data;
  output [15:0] dataOut;
  input clk, reset, write;
  wire   n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n100, n101;

  DFFR_X1 \Reg_reg[15]  ( .D(n53), .CK(clk), .RN(n54), .Q(dataOut[15]), .QN(
        n70) );
  DFFR_X1 \Reg_reg[14]  ( .D(n55), .CK(clk), .RN(n54), .Q(dataOut[14]), .QN(
        n71) );
  DFFR_X1 \Reg_reg[13]  ( .D(n56), .CK(clk), .RN(n54), .Q(dataOut[13]), .QN(
        n72) );
  DFFR_X1 \Reg_reg[12]  ( .D(n57), .CK(clk), .RN(n54), .Q(dataOut[12]), .QN(
        n73) );
  DFFR_X1 \Reg_reg[11]  ( .D(n58), .CK(clk), .RN(n54), .Q(dataOut[11]), .QN(
        n74) );
  DFFR_X1 \Reg_reg[10]  ( .D(n59), .CK(clk), .RN(n54), .Q(dataOut[10]), .QN(
        n75) );
  DFFR_X1 \Reg_reg[9]  ( .D(n60), .CK(clk), .RN(n54), .Q(dataOut[9]), .QN(n76)
         );
  DFFR_X1 \Reg_reg[8]  ( .D(n61), .CK(clk), .RN(n54), .Q(dataOut[8]), .QN(n77)
         );
  DFFR_X1 \Reg_reg[7]  ( .D(n62), .CK(clk), .RN(n54), .Q(dataOut[7]), .QN(n78)
         );
  DFFR_X1 \Reg_reg[6]  ( .D(n63), .CK(clk), .RN(n54), .Q(dataOut[6]), .QN(n79)
         );
  DFFR_X1 \Reg_reg[5]  ( .D(n64), .CK(clk), .RN(n54), .Q(dataOut[5]), .QN(n80)
         );
  DFFR_X1 \Reg_reg[4]  ( .D(n65), .CK(clk), .RN(n54), .Q(dataOut[4]), .QN(n81)
         );
  DFFR_X1 \Reg_reg[3]  ( .D(n66), .CK(clk), .RN(n54), .Q(dataOut[3]), .QN(n82)
         );
  DFFR_X1 \Reg_reg[2]  ( .D(n67), .CK(clk), .RN(n54), .Q(dataOut[2]), .QN(n83)
         );
  DFFR_X1 \Reg_reg[1]  ( .D(n68), .CK(clk), .RN(n54), .Q(dataOut[1]), .QN(n84)
         );
  DFFR_X1 \Reg_reg[0]  ( .D(n69), .CK(clk), .RN(n54), .Q(dataOut[0]), .QN(n85)
         );
  OAI21_X1 U2 ( .B1(n50), .B2(n85), .A(n101), .ZN(n69) );
  NAND2_X1 U3 ( .A1(n52), .A2(data[0]), .ZN(n101) );
  OAI21_X1 U4 ( .B1(n50), .B2(n84), .A(n100), .ZN(n68) );
  NAND2_X1 U5 ( .A1(data[1]), .A2(n52), .ZN(n100) );
  OAI21_X1 U6 ( .B1(n50), .B2(n83), .A(n99), .ZN(n67) );
  NAND2_X1 U7 ( .A1(data[2]), .A2(n52), .ZN(n99) );
  OAI21_X1 U8 ( .B1(n50), .B2(n82), .A(n98), .ZN(n66) );
  NAND2_X1 U9 ( .A1(data[3]), .A2(n52), .ZN(n98) );
  OAI21_X1 U10 ( .B1(n50), .B2(n81), .A(n97), .ZN(n65) );
  NAND2_X1 U11 ( .A1(data[4]), .A2(n52), .ZN(n97) );
  OAI21_X1 U12 ( .B1(n50), .B2(n80), .A(n96), .ZN(n64) );
  NAND2_X1 U13 ( .A1(data[5]), .A2(n52), .ZN(n96) );
  OAI21_X1 U14 ( .B1(n50), .B2(n79), .A(n95), .ZN(n63) );
  NAND2_X1 U15 ( .A1(data[6]), .A2(n52), .ZN(n95) );
  OAI21_X1 U16 ( .B1(n51), .B2(n78), .A(n94), .ZN(n62) );
  NAND2_X1 U17 ( .A1(data[7]), .A2(n52), .ZN(n94) );
  OAI21_X1 U18 ( .B1(n51), .B2(n77), .A(n93), .ZN(n61) );
  NAND2_X1 U19 ( .A1(data[8]), .A2(n51), .ZN(n93) );
  OAI21_X1 U20 ( .B1(n51), .B2(n76), .A(n92), .ZN(n60) );
  NAND2_X1 U21 ( .A1(data[9]), .A2(n51), .ZN(n92) );
  OAI21_X1 U22 ( .B1(n50), .B2(n75), .A(n91), .ZN(n59) );
  NAND2_X1 U23 ( .A1(data[10]), .A2(n51), .ZN(n91) );
  OAI21_X1 U24 ( .B1(n51), .B2(n74), .A(n90), .ZN(n58) );
  NAND2_X1 U25 ( .A1(data[11]), .A2(n51), .ZN(n90) );
  OAI21_X1 U26 ( .B1(n50), .B2(n73), .A(n89), .ZN(n57) );
  NAND2_X1 U27 ( .A1(data[12]), .A2(n51), .ZN(n89) );
  OAI21_X1 U28 ( .B1(n50), .B2(n72), .A(n88), .ZN(n56) );
  NAND2_X1 U29 ( .A1(data[13]), .A2(n51), .ZN(n88) );
  OAI21_X1 U30 ( .B1(n50), .B2(n71), .A(n87), .ZN(n55) );
  NAND2_X1 U31 ( .A1(data[14]), .A2(n51), .ZN(n87) );
  INV_X1 U32 ( .A(reset), .ZN(n54) );
  OAI21_X1 U33 ( .B1(n50), .B2(n70), .A(n86), .ZN(n53) );
  NAND2_X1 U34 ( .A1(data[15]), .A2(n51), .ZN(n86) );
  CLKBUF_X3 U35 ( .A(write), .Z(n50) );
  CLKBUF_X3 U36 ( .A(write), .Z(n51) );
  CLKBUF_X3 U37 ( .A(write), .Z(n52) );
endmodule


module SingleReg_7 ( data, clk, reset, write, dataOut );
  input [15:0] data;
  output [15:0] dataOut;
  input clk, reset, write;
  wire   n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n100, n101;

  DFFR_X1 \Reg_reg[15]  ( .D(n53), .CK(clk), .RN(n54), .Q(dataOut[15]), .QN(
        n70) );
  DFFR_X1 \Reg_reg[14]  ( .D(n55), .CK(clk), .RN(n54), .Q(dataOut[14]), .QN(
        n71) );
  DFFR_X1 \Reg_reg[13]  ( .D(n56), .CK(clk), .RN(n54), .Q(dataOut[13]), .QN(
        n72) );
  DFFR_X1 \Reg_reg[12]  ( .D(n57), .CK(clk), .RN(n54), .Q(dataOut[12]), .QN(
        n73) );
  DFFR_X1 \Reg_reg[11]  ( .D(n58), .CK(clk), .RN(n54), .Q(dataOut[11]), .QN(
        n74) );
  DFFR_X1 \Reg_reg[10]  ( .D(n59), .CK(clk), .RN(n54), .Q(dataOut[10]), .QN(
        n75) );
  DFFR_X1 \Reg_reg[9]  ( .D(n60), .CK(clk), .RN(n54), .Q(dataOut[9]), .QN(n76)
         );
  DFFR_X1 \Reg_reg[8]  ( .D(n61), .CK(clk), .RN(n54), .Q(dataOut[8]), .QN(n77)
         );
  DFFR_X1 \Reg_reg[7]  ( .D(n62), .CK(clk), .RN(n54), .Q(dataOut[7]), .QN(n78)
         );
  DFFR_X1 \Reg_reg[6]  ( .D(n63), .CK(clk), .RN(n54), .Q(dataOut[6]), .QN(n79)
         );
  DFFR_X1 \Reg_reg[5]  ( .D(n64), .CK(clk), .RN(n54), .Q(dataOut[5]), .QN(n80)
         );
  DFFR_X1 \Reg_reg[4]  ( .D(n65), .CK(clk), .RN(n54), .Q(dataOut[4]), .QN(n81)
         );
  DFFR_X1 \Reg_reg[3]  ( .D(n66), .CK(clk), .RN(n54), .Q(dataOut[3]), .QN(n82)
         );
  DFFR_X1 \Reg_reg[2]  ( .D(n67), .CK(clk), .RN(n54), .Q(dataOut[2]), .QN(n83)
         );
  DFFR_X1 \Reg_reg[1]  ( .D(n68), .CK(clk), .RN(n54), .Q(dataOut[1]), .QN(n84)
         );
  DFFR_X1 \Reg_reg[0]  ( .D(n69), .CK(clk), .RN(n54), .Q(dataOut[0]), .QN(n85)
         );
  OAI21_X1 U2 ( .B1(n50), .B2(n85), .A(n101), .ZN(n69) );
  NAND2_X1 U3 ( .A1(n52), .A2(data[0]), .ZN(n101) );
  OAI21_X1 U4 ( .B1(n50), .B2(n84), .A(n100), .ZN(n68) );
  NAND2_X1 U5 ( .A1(data[1]), .A2(n52), .ZN(n100) );
  OAI21_X1 U6 ( .B1(n50), .B2(n83), .A(n99), .ZN(n67) );
  NAND2_X1 U7 ( .A1(data[2]), .A2(n52), .ZN(n99) );
  OAI21_X1 U8 ( .B1(n50), .B2(n82), .A(n98), .ZN(n66) );
  NAND2_X1 U9 ( .A1(data[3]), .A2(n52), .ZN(n98) );
  OAI21_X1 U10 ( .B1(n50), .B2(n81), .A(n97), .ZN(n65) );
  NAND2_X1 U11 ( .A1(data[4]), .A2(n52), .ZN(n97) );
  OAI21_X1 U12 ( .B1(n50), .B2(n80), .A(n96), .ZN(n64) );
  NAND2_X1 U13 ( .A1(data[5]), .A2(n52), .ZN(n96) );
  OAI21_X1 U14 ( .B1(n50), .B2(n79), .A(n95), .ZN(n63) );
  NAND2_X1 U15 ( .A1(data[6]), .A2(n52), .ZN(n95) );
  OAI21_X1 U16 ( .B1(n51), .B2(n78), .A(n94), .ZN(n62) );
  NAND2_X1 U17 ( .A1(data[7]), .A2(n52), .ZN(n94) );
  OAI21_X1 U18 ( .B1(n51), .B2(n77), .A(n93), .ZN(n61) );
  NAND2_X1 U19 ( .A1(data[8]), .A2(n51), .ZN(n93) );
  OAI21_X1 U20 ( .B1(n51), .B2(n76), .A(n92), .ZN(n60) );
  NAND2_X1 U21 ( .A1(data[9]), .A2(n51), .ZN(n92) );
  OAI21_X1 U22 ( .B1(n50), .B2(n75), .A(n91), .ZN(n59) );
  NAND2_X1 U23 ( .A1(data[10]), .A2(n51), .ZN(n91) );
  OAI21_X1 U24 ( .B1(n51), .B2(n74), .A(n90), .ZN(n58) );
  NAND2_X1 U25 ( .A1(data[11]), .A2(n51), .ZN(n90) );
  OAI21_X1 U26 ( .B1(n50), .B2(n73), .A(n89), .ZN(n57) );
  NAND2_X1 U27 ( .A1(data[12]), .A2(n51), .ZN(n89) );
  OAI21_X1 U28 ( .B1(n50), .B2(n72), .A(n88), .ZN(n56) );
  NAND2_X1 U29 ( .A1(data[13]), .A2(n51), .ZN(n88) );
  OAI21_X1 U30 ( .B1(n50), .B2(n71), .A(n87), .ZN(n55) );
  NAND2_X1 U31 ( .A1(data[14]), .A2(n51), .ZN(n87) );
  INV_X1 U32 ( .A(reset), .ZN(n54) );
  OAI21_X1 U33 ( .B1(n50), .B2(n70), .A(n86), .ZN(n53) );
  NAND2_X1 U34 ( .A1(data[15]), .A2(n51), .ZN(n86) );
  CLKBUF_X3 U35 ( .A(write), .Z(n50) );
  CLKBUF_X3 U36 ( .A(write), .Z(n51) );
  CLKBUF_X3 U37 ( .A(write), .Z(n52) );
endmodule


module SingleReg_6 ( data, clk, reset, write, dataOut );
  input [15:0] data;
  output [15:0] dataOut;
  input clk, reset, write;
  wire   n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n100, n101;

  DFFR_X1 \Reg_reg[15]  ( .D(n53), .CK(clk), .RN(n54), .Q(dataOut[15]), .QN(
        n70) );
  DFFR_X1 \Reg_reg[14]  ( .D(n55), .CK(clk), .RN(n54), .Q(dataOut[14]), .QN(
        n71) );
  DFFR_X1 \Reg_reg[13]  ( .D(n56), .CK(clk), .RN(n54), .Q(dataOut[13]), .QN(
        n72) );
  DFFR_X1 \Reg_reg[12]  ( .D(n57), .CK(clk), .RN(n54), .Q(dataOut[12]), .QN(
        n73) );
  DFFR_X1 \Reg_reg[11]  ( .D(n58), .CK(clk), .RN(n54), .Q(dataOut[11]), .QN(
        n74) );
  DFFR_X1 \Reg_reg[10]  ( .D(n59), .CK(clk), .RN(n54), .Q(dataOut[10]), .QN(
        n75) );
  DFFR_X1 \Reg_reg[9]  ( .D(n60), .CK(clk), .RN(n54), .Q(dataOut[9]), .QN(n76)
         );
  DFFR_X1 \Reg_reg[8]  ( .D(n61), .CK(clk), .RN(n54), .Q(dataOut[8]), .QN(n77)
         );
  DFFR_X1 \Reg_reg[7]  ( .D(n62), .CK(clk), .RN(n54), .Q(dataOut[7]), .QN(n78)
         );
  DFFR_X1 \Reg_reg[6]  ( .D(n63), .CK(clk), .RN(n54), .Q(dataOut[6]), .QN(n79)
         );
  DFFR_X1 \Reg_reg[5]  ( .D(n64), .CK(clk), .RN(n54), .Q(dataOut[5]), .QN(n80)
         );
  DFFR_X1 \Reg_reg[4]  ( .D(n65), .CK(clk), .RN(n54), .Q(dataOut[4]), .QN(n81)
         );
  DFFR_X1 \Reg_reg[3]  ( .D(n66), .CK(clk), .RN(n54), .Q(dataOut[3]), .QN(n82)
         );
  DFFR_X1 \Reg_reg[2]  ( .D(n67), .CK(clk), .RN(n54), .Q(dataOut[2]), .QN(n83)
         );
  DFFR_X1 \Reg_reg[1]  ( .D(n68), .CK(clk), .RN(n54), .Q(dataOut[1]), .QN(n84)
         );
  DFFR_X1 \Reg_reg[0]  ( .D(n69), .CK(clk), .RN(n54), .Q(dataOut[0]), .QN(n85)
         );
  OAI21_X1 U2 ( .B1(n50), .B2(n85), .A(n101), .ZN(n69) );
  NAND2_X1 U3 ( .A1(n52), .A2(data[0]), .ZN(n101) );
  OAI21_X1 U4 ( .B1(n50), .B2(n84), .A(n100), .ZN(n68) );
  NAND2_X1 U5 ( .A1(data[1]), .A2(n52), .ZN(n100) );
  OAI21_X1 U6 ( .B1(n50), .B2(n83), .A(n99), .ZN(n67) );
  NAND2_X1 U7 ( .A1(data[2]), .A2(n52), .ZN(n99) );
  OAI21_X1 U8 ( .B1(n50), .B2(n82), .A(n98), .ZN(n66) );
  NAND2_X1 U9 ( .A1(data[3]), .A2(n52), .ZN(n98) );
  OAI21_X1 U10 ( .B1(n50), .B2(n81), .A(n97), .ZN(n65) );
  NAND2_X1 U11 ( .A1(data[4]), .A2(n52), .ZN(n97) );
  OAI21_X1 U12 ( .B1(n50), .B2(n80), .A(n96), .ZN(n64) );
  NAND2_X1 U13 ( .A1(data[5]), .A2(n52), .ZN(n96) );
  OAI21_X1 U14 ( .B1(n50), .B2(n79), .A(n95), .ZN(n63) );
  NAND2_X1 U15 ( .A1(data[6]), .A2(n52), .ZN(n95) );
  OAI21_X1 U16 ( .B1(n51), .B2(n78), .A(n94), .ZN(n62) );
  NAND2_X1 U17 ( .A1(data[7]), .A2(n52), .ZN(n94) );
  OAI21_X1 U18 ( .B1(n51), .B2(n77), .A(n93), .ZN(n61) );
  NAND2_X1 U19 ( .A1(data[8]), .A2(n51), .ZN(n93) );
  OAI21_X1 U20 ( .B1(n51), .B2(n76), .A(n92), .ZN(n60) );
  NAND2_X1 U21 ( .A1(data[9]), .A2(n51), .ZN(n92) );
  OAI21_X1 U22 ( .B1(n50), .B2(n75), .A(n91), .ZN(n59) );
  NAND2_X1 U23 ( .A1(data[10]), .A2(n51), .ZN(n91) );
  OAI21_X1 U24 ( .B1(n51), .B2(n74), .A(n90), .ZN(n58) );
  NAND2_X1 U25 ( .A1(data[11]), .A2(n51), .ZN(n90) );
  OAI21_X1 U26 ( .B1(n50), .B2(n73), .A(n89), .ZN(n57) );
  NAND2_X1 U27 ( .A1(data[12]), .A2(n51), .ZN(n89) );
  OAI21_X1 U28 ( .B1(n50), .B2(n72), .A(n88), .ZN(n56) );
  NAND2_X1 U29 ( .A1(data[13]), .A2(n51), .ZN(n88) );
  OAI21_X1 U30 ( .B1(n50), .B2(n71), .A(n87), .ZN(n55) );
  NAND2_X1 U31 ( .A1(data[14]), .A2(n51), .ZN(n87) );
  INV_X1 U32 ( .A(reset), .ZN(n54) );
  OAI21_X1 U33 ( .B1(n50), .B2(n70), .A(n86), .ZN(n53) );
  NAND2_X1 U34 ( .A1(data[15]), .A2(n51), .ZN(n86) );
  CLKBUF_X3 U35 ( .A(write), .Z(n50) );
  CLKBUF_X3 U36 ( .A(write), .Z(n51) );
  CLKBUF_X3 U37 ( .A(write), .Z(n52) );
endmodule


module SingleReg_5 ( data, clk, reset, write, dataOut );
  input [15:0] data;
  output [15:0] dataOut;
  input clk, reset, write;
  wire   n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n100, n101;

  DFFR_X1 \Reg_reg[15]  ( .D(n53), .CK(clk), .RN(n54), .Q(dataOut[15]), .QN(
        n70) );
  DFFR_X1 \Reg_reg[14]  ( .D(n55), .CK(clk), .RN(n54), .Q(dataOut[14]), .QN(
        n71) );
  DFFR_X1 \Reg_reg[13]  ( .D(n56), .CK(clk), .RN(n54), .Q(dataOut[13]), .QN(
        n72) );
  DFFR_X1 \Reg_reg[12]  ( .D(n57), .CK(clk), .RN(n54), .Q(dataOut[12]), .QN(
        n73) );
  DFFR_X1 \Reg_reg[11]  ( .D(n58), .CK(clk), .RN(n54), .Q(dataOut[11]), .QN(
        n74) );
  DFFR_X1 \Reg_reg[10]  ( .D(n59), .CK(clk), .RN(n54), .Q(dataOut[10]), .QN(
        n75) );
  DFFR_X1 \Reg_reg[9]  ( .D(n60), .CK(clk), .RN(n54), .Q(dataOut[9]), .QN(n76)
         );
  DFFR_X1 \Reg_reg[8]  ( .D(n61), .CK(clk), .RN(n54), .Q(dataOut[8]), .QN(n77)
         );
  DFFR_X1 \Reg_reg[7]  ( .D(n62), .CK(clk), .RN(n54), .Q(dataOut[7]), .QN(n78)
         );
  DFFR_X1 \Reg_reg[6]  ( .D(n63), .CK(clk), .RN(n54), .Q(dataOut[6]), .QN(n79)
         );
  DFFR_X1 \Reg_reg[5]  ( .D(n64), .CK(clk), .RN(n54), .Q(dataOut[5]), .QN(n80)
         );
  DFFR_X1 \Reg_reg[4]  ( .D(n65), .CK(clk), .RN(n54), .Q(dataOut[4]), .QN(n81)
         );
  DFFR_X1 \Reg_reg[3]  ( .D(n66), .CK(clk), .RN(n54), .Q(dataOut[3]), .QN(n82)
         );
  DFFR_X1 \Reg_reg[2]  ( .D(n67), .CK(clk), .RN(n54), .Q(dataOut[2]), .QN(n83)
         );
  DFFR_X1 \Reg_reg[1]  ( .D(n68), .CK(clk), .RN(n54), .Q(dataOut[1]), .QN(n84)
         );
  DFFR_X1 \Reg_reg[0]  ( .D(n69), .CK(clk), .RN(n54), .Q(dataOut[0]), .QN(n85)
         );
  OAI21_X1 U2 ( .B1(n50), .B2(n85), .A(n101), .ZN(n69) );
  NAND2_X1 U3 ( .A1(n52), .A2(data[0]), .ZN(n101) );
  OAI21_X1 U4 ( .B1(n50), .B2(n84), .A(n100), .ZN(n68) );
  NAND2_X1 U5 ( .A1(data[1]), .A2(n52), .ZN(n100) );
  OAI21_X1 U6 ( .B1(n50), .B2(n83), .A(n99), .ZN(n67) );
  NAND2_X1 U7 ( .A1(data[2]), .A2(n52), .ZN(n99) );
  OAI21_X1 U8 ( .B1(n50), .B2(n82), .A(n98), .ZN(n66) );
  NAND2_X1 U9 ( .A1(data[3]), .A2(n52), .ZN(n98) );
  OAI21_X1 U10 ( .B1(n50), .B2(n81), .A(n97), .ZN(n65) );
  NAND2_X1 U11 ( .A1(data[4]), .A2(n52), .ZN(n97) );
  OAI21_X1 U12 ( .B1(n50), .B2(n80), .A(n96), .ZN(n64) );
  NAND2_X1 U13 ( .A1(data[5]), .A2(n52), .ZN(n96) );
  OAI21_X1 U14 ( .B1(n50), .B2(n79), .A(n95), .ZN(n63) );
  NAND2_X1 U15 ( .A1(data[6]), .A2(n52), .ZN(n95) );
  OAI21_X1 U16 ( .B1(n51), .B2(n78), .A(n94), .ZN(n62) );
  NAND2_X1 U17 ( .A1(data[7]), .A2(n52), .ZN(n94) );
  OAI21_X1 U18 ( .B1(n51), .B2(n77), .A(n93), .ZN(n61) );
  NAND2_X1 U19 ( .A1(data[8]), .A2(n51), .ZN(n93) );
  OAI21_X1 U20 ( .B1(n51), .B2(n76), .A(n92), .ZN(n60) );
  NAND2_X1 U21 ( .A1(data[9]), .A2(n51), .ZN(n92) );
  OAI21_X1 U22 ( .B1(n50), .B2(n75), .A(n91), .ZN(n59) );
  NAND2_X1 U23 ( .A1(data[10]), .A2(n51), .ZN(n91) );
  OAI21_X1 U24 ( .B1(n51), .B2(n74), .A(n90), .ZN(n58) );
  NAND2_X1 U25 ( .A1(data[11]), .A2(n51), .ZN(n90) );
  OAI21_X1 U26 ( .B1(n50), .B2(n73), .A(n89), .ZN(n57) );
  NAND2_X1 U27 ( .A1(data[12]), .A2(n51), .ZN(n89) );
  OAI21_X1 U28 ( .B1(n50), .B2(n72), .A(n88), .ZN(n56) );
  NAND2_X1 U29 ( .A1(data[13]), .A2(n51), .ZN(n88) );
  OAI21_X1 U30 ( .B1(n50), .B2(n71), .A(n87), .ZN(n55) );
  NAND2_X1 U31 ( .A1(data[14]), .A2(n51), .ZN(n87) );
  INV_X1 U32 ( .A(reset), .ZN(n54) );
  OAI21_X1 U33 ( .B1(n50), .B2(n70), .A(n86), .ZN(n53) );
  NAND2_X1 U34 ( .A1(data[15]), .A2(n51), .ZN(n86) );
  CLKBUF_X3 U35 ( .A(write), .Z(n50) );
  CLKBUF_X3 U36 ( .A(write), .Z(n51) );
  CLKBUF_X3 U37 ( .A(write), .Z(n52) );
endmodule


module SingleReg_4 ( data, clk, reset, write, dataOut );
  input [15:0] data;
  output [15:0] dataOut;
  input clk, reset, write;
  wire   n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n100, n101;

  DFFR_X1 \Reg_reg[15]  ( .D(n53), .CK(clk), .RN(n54), .Q(dataOut[15]), .QN(
        n70) );
  DFFR_X1 \Reg_reg[14]  ( .D(n55), .CK(clk), .RN(n54), .Q(dataOut[14]), .QN(
        n71) );
  DFFR_X1 \Reg_reg[13]  ( .D(n56), .CK(clk), .RN(n54), .Q(dataOut[13]), .QN(
        n72) );
  DFFR_X1 \Reg_reg[12]  ( .D(n57), .CK(clk), .RN(n54), .Q(dataOut[12]), .QN(
        n73) );
  DFFR_X1 \Reg_reg[11]  ( .D(n58), .CK(clk), .RN(n54), .Q(dataOut[11]), .QN(
        n74) );
  DFFR_X1 \Reg_reg[10]  ( .D(n59), .CK(clk), .RN(n54), .Q(dataOut[10]), .QN(
        n75) );
  DFFR_X1 \Reg_reg[9]  ( .D(n60), .CK(clk), .RN(n54), .Q(dataOut[9]), .QN(n76)
         );
  DFFR_X1 \Reg_reg[8]  ( .D(n61), .CK(clk), .RN(n54), .Q(dataOut[8]), .QN(n77)
         );
  DFFR_X1 \Reg_reg[7]  ( .D(n62), .CK(clk), .RN(n54), .Q(dataOut[7]), .QN(n78)
         );
  DFFR_X1 \Reg_reg[6]  ( .D(n63), .CK(clk), .RN(n54), .Q(dataOut[6]), .QN(n79)
         );
  DFFR_X1 \Reg_reg[5]  ( .D(n64), .CK(clk), .RN(n54), .Q(dataOut[5]), .QN(n80)
         );
  DFFR_X1 \Reg_reg[4]  ( .D(n65), .CK(clk), .RN(n54), .Q(dataOut[4]), .QN(n81)
         );
  DFFR_X1 \Reg_reg[3]  ( .D(n66), .CK(clk), .RN(n54), .Q(dataOut[3]), .QN(n82)
         );
  DFFR_X1 \Reg_reg[2]  ( .D(n67), .CK(clk), .RN(n54), .Q(dataOut[2]), .QN(n83)
         );
  DFFR_X1 \Reg_reg[1]  ( .D(n68), .CK(clk), .RN(n54), .Q(dataOut[1]), .QN(n84)
         );
  DFFR_X1 \Reg_reg[0]  ( .D(n69), .CK(clk), .RN(n54), .Q(dataOut[0]), .QN(n85)
         );
  OAI21_X1 U2 ( .B1(n50), .B2(n85), .A(n101), .ZN(n69) );
  NAND2_X1 U3 ( .A1(n52), .A2(data[0]), .ZN(n101) );
  OAI21_X1 U4 ( .B1(n50), .B2(n84), .A(n100), .ZN(n68) );
  NAND2_X1 U5 ( .A1(data[1]), .A2(n52), .ZN(n100) );
  OAI21_X1 U6 ( .B1(n50), .B2(n83), .A(n99), .ZN(n67) );
  NAND2_X1 U7 ( .A1(data[2]), .A2(n52), .ZN(n99) );
  OAI21_X1 U8 ( .B1(n50), .B2(n82), .A(n98), .ZN(n66) );
  NAND2_X1 U9 ( .A1(data[3]), .A2(n52), .ZN(n98) );
  OAI21_X1 U10 ( .B1(n50), .B2(n81), .A(n97), .ZN(n65) );
  NAND2_X1 U11 ( .A1(data[4]), .A2(n52), .ZN(n97) );
  OAI21_X1 U12 ( .B1(n50), .B2(n80), .A(n96), .ZN(n64) );
  NAND2_X1 U13 ( .A1(data[5]), .A2(n52), .ZN(n96) );
  OAI21_X1 U14 ( .B1(n50), .B2(n79), .A(n95), .ZN(n63) );
  NAND2_X1 U15 ( .A1(data[6]), .A2(n52), .ZN(n95) );
  OAI21_X1 U16 ( .B1(n51), .B2(n78), .A(n94), .ZN(n62) );
  NAND2_X1 U17 ( .A1(data[7]), .A2(n52), .ZN(n94) );
  OAI21_X1 U18 ( .B1(n51), .B2(n77), .A(n93), .ZN(n61) );
  NAND2_X1 U19 ( .A1(data[8]), .A2(n51), .ZN(n93) );
  OAI21_X1 U20 ( .B1(n51), .B2(n76), .A(n92), .ZN(n60) );
  NAND2_X1 U21 ( .A1(data[9]), .A2(n51), .ZN(n92) );
  OAI21_X1 U22 ( .B1(n50), .B2(n75), .A(n91), .ZN(n59) );
  NAND2_X1 U23 ( .A1(data[10]), .A2(n51), .ZN(n91) );
  OAI21_X1 U24 ( .B1(n51), .B2(n74), .A(n90), .ZN(n58) );
  NAND2_X1 U25 ( .A1(data[11]), .A2(n51), .ZN(n90) );
  OAI21_X1 U26 ( .B1(n50), .B2(n73), .A(n89), .ZN(n57) );
  NAND2_X1 U27 ( .A1(data[12]), .A2(n51), .ZN(n89) );
  OAI21_X1 U28 ( .B1(n50), .B2(n72), .A(n88), .ZN(n56) );
  NAND2_X1 U29 ( .A1(data[13]), .A2(n51), .ZN(n88) );
  OAI21_X1 U30 ( .B1(n50), .B2(n71), .A(n87), .ZN(n55) );
  NAND2_X1 U31 ( .A1(data[14]), .A2(n51), .ZN(n87) );
  INV_X1 U32 ( .A(reset), .ZN(n54) );
  OAI21_X1 U33 ( .B1(n50), .B2(n70), .A(n86), .ZN(n53) );
  NAND2_X1 U34 ( .A1(data[15]), .A2(n51), .ZN(n86) );
  CLKBUF_X3 U35 ( .A(write), .Z(n50) );
  CLKBUF_X3 U36 ( .A(write), .Z(n51) );
  CLKBUF_X3 U37 ( .A(write), .Z(n52) );
endmodule


module SingleReg_3 ( data, clk, reset, write, dataOut );
  input [15:0] data;
  output [15:0] dataOut;
  input clk, reset, write;
  wire   n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n100, n101;

  DFFR_X1 \Reg_reg[15]  ( .D(n53), .CK(clk), .RN(n54), .Q(dataOut[15]), .QN(
        n70) );
  DFFR_X1 \Reg_reg[14]  ( .D(n55), .CK(clk), .RN(n54), .Q(dataOut[14]), .QN(
        n71) );
  DFFR_X1 \Reg_reg[13]  ( .D(n56), .CK(clk), .RN(n54), .Q(dataOut[13]), .QN(
        n72) );
  DFFR_X1 \Reg_reg[12]  ( .D(n57), .CK(clk), .RN(n54), .Q(dataOut[12]), .QN(
        n73) );
  DFFR_X1 \Reg_reg[11]  ( .D(n58), .CK(clk), .RN(n54), .Q(dataOut[11]), .QN(
        n74) );
  DFFR_X1 \Reg_reg[10]  ( .D(n59), .CK(clk), .RN(n54), .Q(dataOut[10]), .QN(
        n75) );
  DFFR_X1 \Reg_reg[9]  ( .D(n60), .CK(clk), .RN(n54), .Q(dataOut[9]), .QN(n76)
         );
  DFFR_X1 \Reg_reg[8]  ( .D(n61), .CK(clk), .RN(n54), .Q(dataOut[8]), .QN(n77)
         );
  DFFR_X1 \Reg_reg[7]  ( .D(n62), .CK(clk), .RN(n54), .Q(dataOut[7]), .QN(n78)
         );
  DFFR_X1 \Reg_reg[6]  ( .D(n63), .CK(clk), .RN(n54), .Q(dataOut[6]), .QN(n79)
         );
  DFFR_X1 \Reg_reg[5]  ( .D(n64), .CK(clk), .RN(n54), .Q(dataOut[5]), .QN(n80)
         );
  DFFR_X1 \Reg_reg[4]  ( .D(n65), .CK(clk), .RN(n54), .Q(dataOut[4]), .QN(n81)
         );
  DFFR_X1 \Reg_reg[3]  ( .D(n66), .CK(clk), .RN(n54), .Q(dataOut[3]), .QN(n82)
         );
  DFFR_X1 \Reg_reg[2]  ( .D(n67), .CK(clk), .RN(n54), .Q(dataOut[2]), .QN(n83)
         );
  DFFR_X1 \Reg_reg[1]  ( .D(n68), .CK(clk), .RN(n54), .Q(dataOut[1]), .QN(n84)
         );
  DFFR_X1 \Reg_reg[0]  ( .D(n69), .CK(clk), .RN(n54), .Q(dataOut[0]), .QN(n85)
         );
  OAI21_X1 U2 ( .B1(n50), .B2(n85), .A(n101), .ZN(n69) );
  NAND2_X1 U3 ( .A1(n52), .A2(data[0]), .ZN(n101) );
  OAI21_X1 U4 ( .B1(n50), .B2(n84), .A(n100), .ZN(n68) );
  NAND2_X1 U5 ( .A1(data[1]), .A2(n52), .ZN(n100) );
  OAI21_X1 U6 ( .B1(n50), .B2(n83), .A(n99), .ZN(n67) );
  NAND2_X1 U7 ( .A1(data[2]), .A2(n52), .ZN(n99) );
  OAI21_X1 U8 ( .B1(n50), .B2(n82), .A(n98), .ZN(n66) );
  NAND2_X1 U9 ( .A1(data[3]), .A2(n52), .ZN(n98) );
  OAI21_X1 U10 ( .B1(n50), .B2(n81), .A(n97), .ZN(n65) );
  NAND2_X1 U11 ( .A1(data[4]), .A2(n52), .ZN(n97) );
  OAI21_X1 U12 ( .B1(n50), .B2(n80), .A(n96), .ZN(n64) );
  NAND2_X1 U13 ( .A1(data[5]), .A2(n52), .ZN(n96) );
  OAI21_X1 U14 ( .B1(n50), .B2(n79), .A(n95), .ZN(n63) );
  NAND2_X1 U15 ( .A1(data[6]), .A2(n52), .ZN(n95) );
  OAI21_X1 U16 ( .B1(n51), .B2(n78), .A(n94), .ZN(n62) );
  NAND2_X1 U17 ( .A1(data[7]), .A2(n52), .ZN(n94) );
  OAI21_X1 U18 ( .B1(n51), .B2(n77), .A(n93), .ZN(n61) );
  NAND2_X1 U19 ( .A1(data[8]), .A2(n51), .ZN(n93) );
  OAI21_X1 U20 ( .B1(n51), .B2(n76), .A(n92), .ZN(n60) );
  NAND2_X1 U21 ( .A1(data[9]), .A2(n51), .ZN(n92) );
  OAI21_X1 U22 ( .B1(n50), .B2(n75), .A(n91), .ZN(n59) );
  NAND2_X1 U23 ( .A1(data[10]), .A2(n51), .ZN(n91) );
  OAI21_X1 U24 ( .B1(n51), .B2(n74), .A(n90), .ZN(n58) );
  NAND2_X1 U25 ( .A1(data[11]), .A2(n51), .ZN(n90) );
  OAI21_X1 U26 ( .B1(n50), .B2(n73), .A(n89), .ZN(n57) );
  NAND2_X1 U27 ( .A1(data[12]), .A2(n51), .ZN(n89) );
  OAI21_X1 U28 ( .B1(n50), .B2(n72), .A(n88), .ZN(n56) );
  NAND2_X1 U29 ( .A1(data[13]), .A2(n51), .ZN(n88) );
  OAI21_X1 U30 ( .B1(n50), .B2(n71), .A(n87), .ZN(n55) );
  NAND2_X1 U31 ( .A1(data[14]), .A2(n51), .ZN(n87) );
  INV_X1 U32 ( .A(reset), .ZN(n54) );
  OAI21_X1 U33 ( .B1(n50), .B2(n70), .A(n86), .ZN(n53) );
  NAND2_X1 U34 ( .A1(data[15]), .A2(n51), .ZN(n86) );
  CLKBUF_X3 U35 ( .A(write), .Z(n50) );
  CLKBUF_X3 U36 ( .A(write), .Z(n51) );
  CLKBUF_X3 U37 ( .A(write), .Z(n52) );
endmodule


module SingleReg_2 ( data, clk, reset, write, dataOut );
  input [15:0] data;
  output [15:0] dataOut;
  input clk, reset, write;
  wire   n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n100, n101;

  DFFR_X1 \Reg_reg[15]  ( .D(n53), .CK(clk), .RN(n54), .Q(dataOut[15]), .QN(
        n70) );
  DFFR_X1 \Reg_reg[14]  ( .D(n55), .CK(clk), .RN(n54), .Q(dataOut[14]), .QN(
        n71) );
  DFFR_X1 \Reg_reg[13]  ( .D(n56), .CK(clk), .RN(n54), .Q(dataOut[13]), .QN(
        n72) );
  DFFR_X1 \Reg_reg[12]  ( .D(n57), .CK(clk), .RN(n54), .Q(dataOut[12]), .QN(
        n73) );
  DFFR_X1 \Reg_reg[11]  ( .D(n58), .CK(clk), .RN(n54), .Q(dataOut[11]), .QN(
        n74) );
  DFFR_X1 \Reg_reg[10]  ( .D(n59), .CK(clk), .RN(n54), .Q(dataOut[10]), .QN(
        n75) );
  DFFR_X1 \Reg_reg[9]  ( .D(n60), .CK(clk), .RN(n54), .Q(dataOut[9]), .QN(n76)
         );
  DFFR_X1 \Reg_reg[8]  ( .D(n61), .CK(clk), .RN(n54), .Q(dataOut[8]), .QN(n77)
         );
  DFFR_X1 \Reg_reg[7]  ( .D(n62), .CK(clk), .RN(n54), .Q(dataOut[7]), .QN(n78)
         );
  DFFR_X1 \Reg_reg[6]  ( .D(n63), .CK(clk), .RN(n54), .Q(dataOut[6]), .QN(n79)
         );
  DFFR_X1 \Reg_reg[5]  ( .D(n64), .CK(clk), .RN(n54), .Q(dataOut[5]), .QN(n80)
         );
  DFFR_X1 \Reg_reg[4]  ( .D(n65), .CK(clk), .RN(n54), .Q(dataOut[4]), .QN(n81)
         );
  DFFR_X1 \Reg_reg[3]  ( .D(n66), .CK(clk), .RN(n54), .Q(dataOut[3]), .QN(n82)
         );
  DFFR_X1 \Reg_reg[2]  ( .D(n67), .CK(clk), .RN(n54), .Q(dataOut[2]), .QN(n83)
         );
  DFFR_X1 \Reg_reg[1]  ( .D(n68), .CK(clk), .RN(n54), .Q(dataOut[1]), .QN(n84)
         );
  DFFR_X1 \Reg_reg[0]  ( .D(n69), .CK(clk), .RN(n54), .Q(dataOut[0]), .QN(n85)
         );
  OAI21_X1 U2 ( .B1(n50), .B2(n85), .A(n101), .ZN(n69) );
  NAND2_X1 U3 ( .A1(n52), .A2(data[0]), .ZN(n101) );
  OAI21_X1 U4 ( .B1(n50), .B2(n84), .A(n100), .ZN(n68) );
  NAND2_X1 U5 ( .A1(data[1]), .A2(n52), .ZN(n100) );
  OAI21_X1 U6 ( .B1(n50), .B2(n83), .A(n99), .ZN(n67) );
  NAND2_X1 U7 ( .A1(data[2]), .A2(n52), .ZN(n99) );
  OAI21_X1 U8 ( .B1(n50), .B2(n82), .A(n98), .ZN(n66) );
  NAND2_X1 U9 ( .A1(data[3]), .A2(n52), .ZN(n98) );
  OAI21_X1 U10 ( .B1(n50), .B2(n81), .A(n97), .ZN(n65) );
  NAND2_X1 U11 ( .A1(data[4]), .A2(n52), .ZN(n97) );
  OAI21_X1 U12 ( .B1(n50), .B2(n80), .A(n96), .ZN(n64) );
  NAND2_X1 U13 ( .A1(data[5]), .A2(n52), .ZN(n96) );
  OAI21_X1 U14 ( .B1(n50), .B2(n79), .A(n95), .ZN(n63) );
  NAND2_X1 U15 ( .A1(data[6]), .A2(n52), .ZN(n95) );
  OAI21_X1 U16 ( .B1(n51), .B2(n78), .A(n94), .ZN(n62) );
  NAND2_X1 U17 ( .A1(data[7]), .A2(n52), .ZN(n94) );
  OAI21_X1 U18 ( .B1(n51), .B2(n77), .A(n93), .ZN(n61) );
  NAND2_X1 U19 ( .A1(data[8]), .A2(n51), .ZN(n93) );
  OAI21_X1 U20 ( .B1(n51), .B2(n76), .A(n92), .ZN(n60) );
  NAND2_X1 U21 ( .A1(data[9]), .A2(n51), .ZN(n92) );
  OAI21_X1 U22 ( .B1(n50), .B2(n75), .A(n91), .ZN(n59) );
  NAND2_X1 U23 ( .A1(data[10]), .A2(n51), .ZN(n91) );
  OAI21_X1 U24 ( .B1(n51), .B2(n74), .A(n90), .ZN(n58) );
  NAND2_X1 U25 ( .A1(data[11]), .A2(n51), .ZN(n90) );
  OAI21_X1 U26 ( .B1(n50), .B2(n73), .A(n89), .ZN(n57) );
  NAND2_X1 U27 ( .A1(data[12]), .A2(n51), .ZN(n89) );
  OAI21_X1 U28 ( .B1(n50), .B2(n72), .A(n88), .ZN(n56) );
  NAND2_X1 U29 ( .A1(data[13]), .A2(n51), .ZN(n88) );
  OAI21_X1 U30 ( .B1(n50), .B2(n71), .A(n87), .ZN(n55) );
  NAND2_X1 U31 ( .A1(data[14]), .A2(n51), .ZN(n87) );
  INV_X1 U32 ( .A(reset), .ZN(n54) );
  OAI21_X1 U33 ( .B1(n50), .B2(n70), .A(n86), .ZN(n53) );
  NAND2_X1 U34 ( .A1(data[15]), .A2(n51), .ZN(n86) );
  CLKBUF_X3 U35 ( .A(write), .Z(n50) );
  CLKBUF_X3 U36 ( .A(write), .Z(n51) );
  CLKBUF_X3 U37 ( .A(write), .Z(n52) );
endmodule


module SingleReg_1 ( data, clk, reset, write, dataOut );
  input [15:0] data;
  output [15:0] dataOut;
  input clk, reset, write;
  wire   n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n100, n101;

  DFFR_X1 \Reg_reg[15]  ( .D(n53), .CK(clk), .RN(n54), .Q(dataOut[15]), .QN(
        n70) );
  DFFR_X1 \Reg_reg[14]  ( .D(n55), .CK(clk), .RN(n54), .Q(dataOut[14]), .QN(
        n71) );
  DFFR_X1 \Reg_reg[13]  ( .D(n56), .CK(clk), .RN(n54), .Q(dataOut[13]), .QN(
        n72) );
  DFFR_X1 \Reg_reg[12]  ( .D(n57), .CK(clk), .RN(n54), .Q(dataOut[12]), .QN(
        n73) );
  DFFR_X1 \Reg_reg[11]  ( .D(n58), .CK(clk), .RN(n54), .Q(dataOut[11]), .QN(
        n74) );
  DFFR_X1 \Reg_reg[10]  ( .D(n59), .CK(clk), .RN(n54), .Q(dataOut[10]), .QN(
        n75) );
  DFFR_X1 \Reg_reg[9]  ( .D(n60), .CK(clk), .RN(n54), .Q(dataOut[9]), .QN(n76)
         );
  DFFR_X1 \Reg_reg[8]  ( .D(n61), .CK(clk), .RN(n54), .Q(dataOut[8]), .QN(n77)
         );
  DFFR_X1 \Reg_reg[7]  ( .D(n62), .CK(clk), .RN(n54), .Q(dataOut[7]), .QN(n78)
         );
  DFFR_X1 \Reg_reg[6]  ( .D(n63), .CK(clk), .RN(n54), .Q(dataOut[6]), .QN(n79)
         );
  DFFR_X1 \Reg_reg[5]  ( .D(n64), .CK(clk), .RN(n54), .Q(dataOut[5]), .QN(n80)
         );
  DFFR_X1 \Reg_reg[4]  ( .D(n65), .CK(clk), .RN(n54), .Q(dataOut[4]), .QN(n81)
         );
  DFFR_X1 \Reg_reg[3]  ( .D(n66), .CK(clk), .RN(n54), .Q(dataOut[3]), .QN(n82)
         );
  DFFR_X1 \Reg_reg[2]  ( .D(n67), .CK(clk), .RN(n54), .Q(dataOut[2]), .QN(n83)
         );
  DFFR_X1 \Reg_reg[1]  ( .D(n68), .CK(clk), .RN(n54), .Q(dataOut[1]), .QN(n84)
         );
  DFFR_X1 \Reg_reg[0]  ( .D(n69), .CK(clk), .RN(n54), .Q(dataOut[0]), .QN(n85)
         );
  OAI21_X1 U2 ( .B1(n50), .B2(n85), .A(n101), .ZN(n69) );
  NAND2_X1 U3 ( .A1(n52), .A2(data[0]), .ZN(n101) );
  OAI21_X1 U4 ( .B1(n50), .B2(n84), .A(n100), .ZN(n68) );
  NAND2_X1 U5 ( .A1(data[1]), .A2(n52), .ZN(n100) );
  OAI21_X1 U6 ( .B1(n50), .B2(n83), .A(n99), .ZN(n67) );
  NAND2_X1 U7 ( .A1(data[2]), .A2(n52), .ZN(n99) );
  OAI21_X1 U8 ( .B1(n50), .B2(n82), .A(n98), .ZN(n66) );
  NAND2_X1 U9 ( .A1(data[3]), .A2(n52), .ZN(n98) );
  OAI21_X1 U10 ( .B1(n50), .B2(n81), .A(n97), .ZN(n65) );
  NAND2_X1 U11 ( .A1(data[4]), .A2(n52), .ZN(n97) );
  OAI21_X1 U12 ( .B1(n50), .B2(n80), .A(n96), .ZN(n64) );
  NAND2_X1 U13 ( .A1(data[5]), .A2(n52), .ZN(n96) );
  OAI21_X1 U14 ( .B1(n50), .B2(n79), .A(n95), .ZN(n63) );
  NAND2_X1 U15 ( .A1(data[6]), .A2(n52), .ZN(n95) );
  OAI21_X1 U16 ( .B1(n51), .B2(n78), .A(n94), .ZN(n62) );
  NAND2_X1 U17 ( .A1(data[7]), .A2(n52), .ZN(n94) );
  OAI21_X1 U18 ( .B1(n51), .B2(n77), .A(n93), .ZN(n61) );
  NAND2_X1 U19 ( .A1(data[8]), .A2(n51), .ZN(n93) );
  OAI21_X1 U20 ( .B1(n51), .B2(n76), .A(n92), .ZN(n60) );
  NAND2_X1 U21 ( .A1(data[9]), .A2(n51), .ZN(n92) );
  OAI21_X1 U22 ( .B1(n50), .B2(n75), .A(n91), .ZN(n59) );
  NAND2_X1 U23 ( .A1(data[10]), .A2(n51), .ZN(n91) );
  OAI21_X1 U24 ( .B1(n51), .B2(n74), .A(n90), .ZN(n58) );
  NAND2_X1 U25 ( .A1(data[11]), .A2(n51), .ZN(n90) );
  OAI21_X1 U26 ( .B1(n50), .B2(n73), .A(n89), .ZN(n57) );
  NAND2_X1 U27 ( .A1(data[12]), .A2(n51), .ZN(n89) );
  OAI21_X1 U28 ( .B1(n50), .B2(n72), .A(n88), .ZN(n56) );
  NAND2_X1 U29 ( .A1(data[13]), .A2(n51), .ZN(n88) );
  OAI21_X1 U30 ( .B1(n50), .B2(n71), .A(n87), .ZN(n55) );
  NAND2_X1 U31 ( .A1(data[14]), .A2(n51), .ZN(n87) );
  INV_X1 U32 ( .A(reset), .ZN(n54) );
  OAI21_X1 U33 ( .B1(n50), .B2(n70), .A(n86), .ZN(n53) );
  NAND2_X1 U34 ( .A1(data[15]), .A2(n51), .ZN(n86) );
  CLKBUF_X3 U35 ( .A(write), .Z(n50) );
  CLKBUF_X3 U36 ( .A(write), .Z(n51) );
  CLKBUF_X3 U37 ( .A(write), .Z(n52) );
endmodule


module SingleReg_0 ( data, clk, reset, write, dataOut );
  input [15:0] data;
  output [15:0] dataOut;
  input clk, reset, write;
  wire   n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n100, n101;

  DFFR_X1 \Reg_reg[15]  ( .D(n53), .CK(clk), .RN(n54), .Q(dataOut[15]), .QN(
        n70) );
  DFFR_X1 \Reg_reg[14]  ( .D(n55), .CK(clk), .RN(n54), .Q(dataOut[14]), .QN(
        n71) );
  DFFR_X1 \Reg_reg[13]  ( .D(n56), .CK(clk), .RN(n54), .Q(dataOut[13]), .QN(
        n72) );
  DFFR_X1 \Reg_reg[12]  ( .D(n57), .CK(clk), .RN(n54), .Q(dataOut[12]), .QN(
        n73) );
  DFFR_X1 \Reg_reg[11]  ( .D(n58), .CK(clk), .RN(n54), .Q(dataOut[11]), .QN(
        n74) );
  DFFR_X1 \Reg_reg[10]  ( .D(n59), .CK(clk), .RN(n54), .Q(dataOut[10]), .QN(
        n75) );
  DFFR_X1 \Reg_reg[9]  ( .D(n60), .CK(clk), .RN(n54), .Q(dataOut[9]), .QN(n76)
         );
  DFFR_X1 \Reg_reg[8]  ( .D(n61), .CK(clk), .RN(n54), .Q(dataOut[8]), .QN(n77)
         );
  DFFR_X1 \Reg_reg[7]  ( .D(n62), .CK(clk), .RN(n54), .Q(dataOut[7]), .QN(n78)
         );
  DFFR_X1 \Reg_reg[6]  ( .D(n63), .CK(clk), .RN(n54), .Q(dataOut[6]), .QN(n79)
         );
  DFFR_X1 \Reg_reg[5]  ( .D(n64), .CK(clk), .RN(n54), .Q(dataOut[5]), .QN(n80)
         );
  DFFR_X1 \Reg_reg[4]  ( .D(n65), .CK(clk), .RN(n54), .Q(dataOut[4]), .QN(n81)
         );
  DFFR_X1 \Reg_reg[3]  ( .D(n66), .CK(clk), .RN(n54), .Q(dataOut[3]), .QN(n82)
         );
  DFFR_X1 \Reg_reg[2]  ( .D(n67), .CK(clk), .RN(n54), .Q(dataOut[2]), .QN(n83)
         );
  DFFR_X1 \Reg_reg[1]  ( .D(n68), .CK(clk), .RN(n54), .Q(dataOut[1]), .QN(n84)
         );
  DFFR_X1 \Reg_reg[0]  ( .D(n69), .CK(clk), .RN(n54), .Q(dataOut[0]), .QN(n85)
         );
  OAI21_X1 U2 ( .B1(n50), .B2(n85), .A(n101), .ZN(n69) );
  NAND2_X1 U3 ( .A1(n52), .A2(data[0]), .ZN(n101) );
  OAI21_X1 U4 ( .B1(n50), .B2(n84), .A(n100), .ZN(n68) );
  NAND2_X1 U5 ( .A1(data[1]), .A2(n52), .ZN(n100) );
  OAI21_X1 U6 ( .B1(n50), .B2(n83), .A(n99), .ZN(n67) );
  NAND2_X1 U7 ( .A1(data[2]), .A2(n52), .ZN(n99) );
  OAI21_X1 U8 ( .B1(n50), .B2(n82), .A(n98), .ZN(n66) );
  NAND2_X1 U9 ( .A1(data[3]), .A2(n52), .ZN(n98) );
  OAI21_X1 U10 ( .B1(n50), .B2(n81), .A(n97), .ZN(n65) );
  NAND2_X1 U11 ( .A1(data[4]), .A2(n52), .ZN(n97) );
  OAI21_X1 U12 ( .B1(n50), .B2(n80), .A(n96), .ZN(n64) );
  NAND2_X1 U13 ( .A1(data[5]), .A2(n52), .ZN(n96) );
  OAI21_X1 U14 ( .B1(n50), .B2(n79), .A(n95), .ZN(n63) );
  NAND2_X1 U15 ( .A1(data[6]), .A2(n52), .ZN(n95) );
  OAI21_X1 U16 ( .B1(n51), .B2(n78), .A(n94), .ZN(n62) );
  NAND2_X1 U17 ( .A1(data[7]), .A2(n52), .ZN(n94) );
  OAI21_X1 U18 ( .B1(n51), .B2(n77), .A(n93), .ZN(n61) );
  NAND2_X1 U19 ( .A1(data[8]), .A2(n51), .ZN(n93) );
  OAI21_X1 U20 ( .B1(n51), .B2(n76), .A(n92), .ZN(n60) );
  NAND2_X1 U21 ( .A1(data[9]), .A2(n51), .ZN(n92) );
  OAI21_X1 U22 ( .B1(n50), .B2(n75), .A(n91), .ZN(n59) );
  NAND2_X1 U23 ( .A1(data[10]), .A2(n51), .ZN(n91) );
  OAI21_X1 U24 ( .B1(n51), .B2(n74), .A(n90), .ZN(n58) );
  NAND2_X1 U25 ( .A1(data[11]), .A2(n51), .ZN(n90) );
  OAI21_X1 U26 ( .B1(n50), .B2(n73), .A(n89), .ZN(n57) );
  NAND2_X1 U27 ( .A1(data[12]), .A2(n51), .ZN(n89) );
  OAI21_X1 U28 ( .B1(n50), .B2(n72), .A(n88), .ZN(n56) );
  NAND2_X1 U29 ( .A1(data[13]), .A2(n51), .ZN(n88) );
  OAI21_X1 U30 ( .B1(n50), .B2(n71), .A(n87), .ZN(n55) );
  NAND2_X1 U31 ( .A1(data[14]), .A2(n51), .ZN(n87) );
  INV_X1 U32 ( .A(reset), .ZN(n54) );
  OAI21_X1 U33 ( .B1(n50), .B2(n70), .A(n86), .ZN(n53) );
  NAND2_X1 U34 ( .A1(data[15]), .A2(n51), .ZN(n86) );
  CLKBUF_X3 U35 ( .A(write), .Z(n50) );
  CLKBUF_X3 U36 ( .A(write), .Z(n51) );
  CLKBUF_X3 U37 ( .A(write), .Z(n52) );
endmodule


module SingleReg_31 ( data, clk, reset, write, dataOut );
  input [15:0] data;
  output [15:0] dataOut;
  input clk, reset, write;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52;

  DFFR_X1 \Reg_reg[15]  ( .D(n49), .CK(clk), .RN(n48), .Q(dataOut[15]), .QN(
        n32) );
  DFFR_X1 \Reg_reg[14]  ( .D(n47), .CK(clk), .RN(n48), .Q(dataOut[14]), .QN(
        n31) );
  DFFR_X1 \Reg_reg[13]  ( .D(n46), .CK(clk), .RN(n48), .Q(dataOut[13]), .QN(
        n30) );
  DFFR_X1 \Reg_reg[12]  ( .D(n45), .CK(clk), .RN(n48), .Q(dataOut[12]), .QN(
        n29) );
  DFFR_X1 \Reg_reg[11]  ( .D(n44), .CK(clk), .RN(n48), .Q(dataOut[11]), .QN(
        n28) );
  DFFR_X1 \Reg_reg[10]  ( .D(n43), .CK(clk), .RN(n48), .Q(dataOut[10]), .QN(
        n27) );
  DFFR_X1 \Reg_reg[9]  ( .D(n42), .CK(clk), .RN(n48), .Q(dataOut[9]), .QN(n26)
         );
  DFFR_X1 \Reg_reg[8]  ( .D(n41), .CK(clk), .RN(n48), .Q(dataOut[8]), .QN(n25)
         );
  DFFR_X1 \Reg_reg[7]  ( .D(n40), .CK(clk), .RN(n48), .Q(dataOut[7]), .QN(n24)
         );
  DFFR_X1 \Reg_reg[6]  ( .D(n39), .CK(clk), .RN(n48), .Q(dataOut[6]), .QN(n23)
         );
  DFFR_X1 \Reg_reg[5]  ( .D(n38), .CK(clk), .RN(n48), .Q(dataOut[5]), .QN(n22)
         );
  DFFR_X1 \Reg_reg[4]  ( .D(n37), .CK(clk), .RN(n48), .Q(dataOut[4]), .QN(n21)
         );
  DFFR_X1 \Reg_reg[3]  ( .D(n36), .CK(clk), .RN(n48), .Q(dataOut[3]), .QN(n20)
         );
  DFFR_X1 \Reg_reg[2]  ( .D(n35), .CK(clk), .RN(n48), .Q(dataOut[2]), .QN(n19)
         );
  DFFR_X1 \Reg_reg[1]  ( .D(n34), .CK(clk), .RN(n48), .Q(dataOut[1]), .QN(n18)
         );
  DFFR_X1 \Reg_reg[0]  ( .D(n33), .CK(clk), .RN(n48), .Q(dataOut[0]), .QN(n17)
         );
  OAI21_X1 U2 ( .B1(n50), .B2(n17), .A(n1), .ZN(n33) );
  NAND2_X1 U3 ( .A1(n52), .A2(data[0]), .ZN(n1) );
  OAI21_X1 U4 ( .B1(n50), .B2(n18), .A(n2), .ZN(n34) );
  NAND2_X1 U5 ( .A1(data[1]), .A2(n52), .ZN(n2) );
  OAI21_X1 U6 ( .B1(n50), .B2(n19), .A(n3), .ZN(n35) );
  NAND2_X1 U7 ( .A1(data[2]), .A2(n52), .ZN(n3) );
  OAI21_X1 U8 ( .B1(n50), .B2(n20), .A(n4), .ZN(n36) );
  NAND2_X1 U9 ( .A1(data[3]), .A2(n52), .ZN(n4) );
  OAI21_X1 U10 ( .B1(n50), .B2(n21), .A(n5), .ZN(n37) );
  NAND2_X1 U11 ( .A1(data[4]), .A2(n52), .ZN(n5) );
  OAI21_X1 U12 ( .B1(n50), .B2(n22), .A(n6), .ZN(n38) );
  NAND2_X1 U13 ( .A1(data[5]), .A2(n52), .ZN(n6) );
  OAI21_X1 U14 ( .B1(n50), .B2(n23), .A(n7), .ZN(n39) );
  NAND2_X1 U15 ( .A1(data[6]), .A2(n52), .ZN(n7) );
  OAI21_X1 U16 ( .B1(n51), .B2(n24), .A(n8), .ZN(n40) );
  NAND2_X1 U17 ( .A1(data[7]), .A2(n52), .ZN(n8) );
  OAI21_X1 U18 ( .B1(n51), .B2(n25), .A(n9), .ZN(n41) );
  NAND2_X1 U19 ( .A1(data[8]), .A2(n51), .ZN(n9) );
  OAI21_X1 U20 ( .B1(n51), .B2(n26), .A(n10), .ZN(n42) );
  NAND2_X1 U21 ( .A1(data[9]), .A2(n51), .ZN(n10) );
  OAI21_X1 U22 ( .B1(n50), .B2(n27), .A(n11), .ZN(n43) );
  NAND2_X1 U23 ( .A1(data[10]), .A2(n51), .ZN(n11) );
  OAI21_X1 U24 ( .B1(n51), .B2(n28), .A(n12), .ZN(n44) );
  NAND2_X1 U25 ( .A1(data[11]), .A2(n51), .ZN(n12) );
  OAI21_X1 U26 ( .B1(n50), .B2(n29), .A(n13), .ZN(n45) );
  NAND2_X1 U27 ( .A1(data[12]), .A2(n51), .ZN(n13) );
  OAI21_X1 U28 ( .B1(n50), .B2(n30), .A(n14), .ZN(n46) );
  NAND2_X1 U29 ( .A1(data[13]), .A2(n51), .ZN(n14) );
  OAI21_X1 U30 ( .B1(n50), .B2(n31), .A(n15), .ZN(n47) );
  NAND2_X1 U31 ( .A1(data[14]), .A2(n51), .ZN(n15) );
  INV_X1 U32 ( .A(reset), .ZN(n48) );
  OAI21_X1 U33 ( .B1(n50), .B2(n32), .A(n16), .ZN(n49) );
  NAND2_X1 U34 ( .A1(data[15]), .A2(n51), .ZN(n16) );
  CLKBUF_X3 U35 ( .A(write), .Z(n50) );
  CLKBUF_X3 U36 ( .A(write), .Z(n51) );
  CLKBUF_X3 U37 ( .A(write), .Z(n52) );
endmodule


module RegFile ( addressA, addressB, dataIn, addressIn, clk, reset, write, 
        outA, outB );
  input [4:0] addressA;
  input [4:0] addressB;
  input [15:0] dataIn;
  input [4:0] addressIn;
  output [15:0] outA;
  output [15:0] outB;
  input clk, reset, write;
  wire   \regOut[0][15] , \regOut[0][14] , \regOut[0][13] , \regOut[0][12] ,
         \regOut[0][11] , \regOut[0][10] , \regOut[0][9] , \regOut[0][8] ,
         \regOut[0][7] , \regOut[0][6] , \regOut[0][5] , \regOut[0][4] ,
         \regOut[0][3] , \regOut[0][2] , \regOut[0][1] , \regOut[0][0] ,
         \regOut[1][15] , \regOut[1][14] , \regOut[1][13] , \regOut[1][12] ,
         \regOut[1][11] , \regOut[1][10] , \regOut[1][9] , \regOut[1][8] ,
         \regOut[1][7] , \regOut[1][6] , \regOut[1][5] , \regOut[1][4] ,
         \regOut[1][3] , \regOut[1][2] , \regOut[1][1] , \regOut[1][0] ,
         \regOut[2][15] , \regOut[2][14] , \regOut[2][13] , \regOut[2][12] ,
         \regOut[2][11] , \regOut[2][10] , \regOut[2][9] , \regOut[2][8] ,
         \regOut[2][7] , \regOut[2][6] , \regOut[2][5] , \regOut[2][4] ,
         \regOut[2][3] , \regOut[2][2] , \regOut[2][1] , \regOut[2][0] ,
         \regOut[3][15] , \regOut[3][14] , \regOut[3][13] , \regOut[3][12] ,
         \regOut[3][11] , \regOut[3][10] , \regOut[3][9] , \regOut[3][8] ,
         \regOut[3][7] , \regOut[3][6] , \regOut[3][5] , \regOut[3][4] ,
         \regOut[3][3] , \regOut[3][2] , \regOut[3][1] , \regOut[3][0] ,
         \regOut[4][15] , \regOut[4][14] , \regOut[4][13] , \regOut[4][12] ,
         \regOut[4][11] , \regOut[4][10] , \regOut[4][9] , \regOut[4][8] ,
         \regOut[4][7] , \regOut[4][6] , \regOut[4][5] , \regOut[4][4] ,
         \regOut[4][3] , \regOut[4][2] , \regOut[4][1] , \regOut[4][0] ,
         \regOut[5][15] , \regOut[5][14] , \regOut[5][13] , \regOut[5][12] ,
         \regOut[5][11] , \regOut[5][10] , \regOut[5][9] , \regOut[5][8] ,
         \regOut[5][7] , \regOut[5][6] , \regOut[5][5] , \regOut[5][4] ,
         \regOut[5][3] , \regOut[5][2] , \regOut[5][1] , \regOut[5][0] ,
         \regOut[6][15] , \regOut[6][14] , \regOut[6][13] , \regOut[6][12] ,
         \regOut[6][11] , \regOut[6][10] , \regOut[6][9] , \regOut[6][8] ,
         \regOut[6][7] , \regOut[6][6] , \regOut[6][5] , \regOut[6][4] ,
         \regOut[6][3] , \regOut[6][2] , \regOut[6][1] , \regOut[6][0] ,
         \regOut[7][15] , \regOut[7][14] , \regOut[7][13] , \regOut[7][12] ,
         \regOut[7][11] , \regOut[7][10] , \regOut[7][9] , \regOut[7][8] ,
         \regOut[7][7] , \regOut[7][6] , \regOut[7][5] , \regOut[7][4] ,
         \regOut[7][3] , \regOut[7][2] , \regOut[7][1] , \regOut[7][0] ,
         \regOut[8][15] , \regOut[8][14] , \regOut[8][13] , \regOut[8][12] ,
         \regOut[8][11] , \regOut[8][10] , \regOut[8][9] , \regOut[8][8] ,
         \regOut[8][7] , \regOut[8][6] , \regOut[8][5] , \regOut[8][4] ,
         \regOut[8][3] , \regOut[8][2] , \regOut[8][1] , \regOut[8][0] ,
         \regOut[9][15] , \regOut[9][14] , \regOut[9][13] , \regOut[9][12] ,
         \regOut[9][11] , \regOut[9][10] , \regOut[9][9] , \regOut[9][8] ,
         \regOut[9][7] , \regOut[9][6] , \regOut[9][5] , \regOut[9][4] ,
         \regOut[9][3] , \regOut[9][2] , \regOut[9][1] , \regOut[9][0] ,
         \regOut[10][15] , \regOut[10][14] , \regOut[10][13] ,
         \regOut[10][12] , \regOut[10][11] , \regOut[10][10] , \regOut[10][9] ,
         \regOut[10][8] , \regOut[10][7] , \regOut[10][6] , \regOut[10][5] ,
         \regOut[10][4] , \regOut[10][3] , \regOut[10][2] , \regOut[10][1] ,
         \regOut[10][0] , \regOut[11][15] , \regOut[11][14] , \regOut[11][13] ,
         \regOut[11][12] , \regOut[11][11] , \regOut[11][10] , \regOut[11][9] ,
         \regOut[11][8] , \regOut[11][7] , \regOut[11][6] , \regOut[11][5] ,
         \regOut[11][4] , \regOut[11][3] , \regOut[11][2] , \regOut[11][1] ,
         \regOut[11][0] , \regOut[12][15] , \regOut[12][14] , \regOut[12][13] ,
         \regOut[12][12] , \regOut[12][11] , \regOut[12][10] , \regOut[12][9] ,
         \regOut[12][8] , \regOut[12][7] , \regOut[12][6] , \regOut[12][5] ,
         \regOut[12][4] , \regOut[12][3] , \regOut[12][2] , \regOut[12][1] ,
         \regOut[12][0] , \regOut[13][15] , \regOut[13][14] , \regOut[13][13] ,
         \regOut[13][12] , \regOut[13][11] , \regOut[13][10] , \regOut[13][9] ,
         \regOut[13][8] , \regOut[13][7] , \regOut[13][6] , \regOut[13][5] ,
         \regOut[13][4] , \regOut[13][3] , \regOut[13][2] , \regOut[13][1] ,
         \regOut[13][0] , \regOut[14][15] , \regOut[14][14] , \regOut[14][13] ,
         \regOut[14][12] , \regOut[14][11] , \regOut[14][10] , \regOut[14][9] ,
         \regOut[14][8] , \regOut[14][7] , \regOut[14][6] , \regOut[14][5] ,
         \regOut[14][4] , \regOut[14][3] , \regOut[14][2] , \regOut[14][1] ,
         \regOut[14][0] , \regOut[15][15] , \regOut[15][14] , \regOut[15][13] ,
         \regOut[15][12] , \regOut[15][11] , \regOut[15][10] , \regOut[15][9] ,
         \regOut[15][8] , \regOut[15][7] , \regOut[15][6] , \regOut[15][5] ,
         \regOut[15][4] , \regOut[15][3] , \regOut[15][2] , \regOut[15][1] ,
         \regOut[15][0] , \regOut[16][15] , \regOut[16][14] , \regOut[16][13] ,
         \regOut[16][12] , \regOut[16][11] , \regOut[16][10] , \regOut[16][9] ,
         \regOut[16][8] , \regOut[16][7] , \regOut[16][6] , \regOut[16][5] ,
         \regOut[16][4] , \regOut[16][3] , \regOut[16][2] , \regOut[16][1] ,
         \regOut[16][0] , \regOut[17][15] , \regOut[17][14] , \regOut[17][13] ,
         \regOut[17][12] , \regOut[17][11] , \regOut[17][10] , \regOut[17][9] ,
         \regOut[17][8] , \regOut[17][7] , \regOut[17][6] , \regOut[17][5] ,
         \regOut[17][4] , \regOut[17][3] , \regOut[17][2] , \regOut[17][1] ,
         \regOut[17][0] , \regOut[18][15] , \regOut[18][14] , \regOut[18][13] ,
         \regOut[18][12] , \regOut[18][11] , \regOut[18][10] , \regOut[18][9] ,
         \regOut[18][8] , \regOut[18][7] , \regOut[18][6] , \regOut[18][5] ,
         \regOut[18][4] , \regOut[18][3] , \regOut[18][2] , \regOut[18][1] ,
         \regOut[18][0] , \regOut[19][15] , \regOut[19][14] , \regOut[19][13] ,
         \regOut[19][12] , \regOut[19][11] , \regOut[19][10] , \regOut[19][9] ,
         \regOut[19][8] , \regOut[19][7] , \regOut[19][6] , \regOut[19][5] ,
         \regOut[19][4] , \regOut[19][3] , \regOut[19][2] , \regOut[19][1] ,
         \regOut[19][0] , \regOut[20][15] , \regOut[20][14] , \regOut[20][13] ,
         \regOut[20][12] , \regOut[20][11] , \regOut[20][10] , \regOut[20][9] ,
         \regOut[20][8] , \regOut[20][7] , \regOut[20][6] , \regOut[20][5] ,
         \regOut[20][4] , \regOut[20][3] , \regOut[20][2] , \regOut[20][1] ,
         \regOut[20][0] , \regOut[21][15] , \regOut[21][14] , \regOut[21][13] ,
         \regOut[21][12] , \regOut[21][11] , \regOut[21][10] , \regOut[21][9] ,
         \regOut[21][8] , \regOut[21][7] , \regOut[21][6] , \regOut[21][5] ,
         \regOut[21][4] , \regOut[21][3] , \regOut[21][2] , \regOut[21][1] ,
         \regOut[21][0] , \regOut[22][15] , \regOut[22][14] , \regOut[22][13] ,
         \regOut[22][12] , \regOut[22][11] , \regOut[22][10] , \regOut[22][9] ,
         \regOut[22][8] , \regOut[22][7] , \regOut[22][6] , \regOut[22][5] ,
         \regOut[22][4] , \regOut[22][3] , \regOut[22][2] , \regOut[22][1] ,
         \regOut[22][0] , \regOut[23][15] , \regOut[23][14] , \regOut[23][13] ,
         \regOut[23][12] , \regOut[23][11] , \regOut[23][10] , \regOut[23][9] ,
         \regOut[23][8] , \regOut[23][7] , \regOut[23][6] , \regOut[23][5] ,
         \regOut[23][4] , \regOut[23][3] , \regOut[23][2] , \regOut[23][1] ,
         \regOut[23][0] , \regOut[24][15] , \regOut[24][14] , \regOut[24][13] ,
         \regOut[24][12] , \regOut[24][11] , \regOut[24][10] , \regOut[24][9] ,
         \regOut[24][8] , \regOut[24][7] , \regOut[24][6] , \regOut[24][5] ,
         \regOut[24][4] , \regOut[24][3] , \regOut[24][2] , \regOut[24][1] ,
         \regOut[24][0] , \regOut[25][15] , \regOut[25][14] , \regOut[25][13] ,
         \regOut[25][12] , \regOut[25][11] , \regOut[25][10] , \regOut[25][9] ,
         \regOut[25][8] , \regOut[25][7] , \regOut[25][6] , \regOut[25][5] ,
         \regOut[25][4] , \regOut[25][3] , \regOut[25][2] , \regOut[25][1] ,
         \regOut[25][0] , \regOut[26][15] , \regOut[26][14] , \regOut[26][13] ,
         \regOut[26][12] , \regOut[26][11] , \regOut[26][10] , \regOut[26][9] ,
         \regOut[26][8] , \regOut[26][7] , \regOut[26][6] , \regOut[26][5] ,
         \regOut[26][4] , \regOut[26][3] , \regOut[26][2] , \regOut[26][1] ,
         \regOut[26][0] , \regOut[27][15] , \regOut[27][14] , \regOut[27][13] ,
         \regOut[27][12] , \regOut[27][11] , \regOut[27][10] , \regOut[27][9] ,
         \regOut[27][8] , \regOut[27][7] , \regOut[27][6] , \regOut[27][5] ,
         \regOut[27][4] , \regOut[27][3] , \regOut[27][2] , \regOut[27][1] ,
         \regOut[27][0] , \regOut[28][15] , \regOut[28][14] , \regOut[28][13] ,
         \regOut[28][12] , \regOut[28][11] , \regOut[28][10] , \regOut[28][9] ,
         \regOut[28][8] , \regOut[28][7] , \regOut[28][6] , \regOut[28][5] ,
         \regOut[28][4] , \regOut[28][3] , \regOut[28][2] , \regOut[28][1] ,
         \regOut[28][0] , \regOut[29][15] , \regOut[29][14] , \regOut[29][13] ,
         \regOut[29][12] , \regOut[29][11] , \regOut[29][10] , \regOut[29][9] ,
         \regOut[29][8] , \regOut[29][7] , \regOut[29][6] , \regOut[29][5] ,
         \regOut[29][4] , \regOut[29][3] , \regOut[29][2] , \regOut[29][1] ,
         \regOut[29][0] , \regOut[30][15] , \regOut[30][14] , \regOut[30][13] ,
         \regOut[30][12] , \regOut[30][11] , \regOut[30][10] , \regOut[30][9] ,
         \regOut[30][8] , \regOut[30][7] , \regOut[30][6] , \regOut[30][5] ,
         \regOut[30][4] , \regOut[30][3] , \regOut[30][2] , \regOut[30][1] ,
         \regOut[30][0] , \regOut[31][15] , \regOut[31][14] , \regOut[31][13] ,
         \regOut[31][12] , \regOut[31][11] , \regOut[31][10] , \regOut[31][9] ,
         \regOut[31][8] , \regOut[31][7] , \regOut[31][6] , \regOut[31][5] ,
         \regOut[31][4] , \regOut[31][3] , \regOut[31][2] , \regOut[31][1] ,
         \regOut[31][0] , \regIn[0][15] , \regIn[0][14] , \regIn[0][13] ,
         \regIn[0][12] , \regIn[0][11] , \regIn[0][10] , \regIn[0][9] ,
         \regIn[0][8] , \regIn[0][7] , \regIn[0][6] , \regIn[0][5] ,
         \regIn[0][4] , \regIn[0][3] , \regIn[0][2] , \regIn[0][1] ,
         \regIn[0][0] , \regIn[1][15] , \regIn[1][14] , \regIn[1][13] ,
         \regIn[1][12] , \regIn[1][11] , \regIn[1][10] , \regIn[1][9] ,
         \regIn[1][8] , \regIn[1][7] , \regIn[1][6] , \regIn[1][5] ,
         \regIn[1][4] , \regIn[1][3] , \regIn[1][2] , \regIn[1][1] ,
         \regIn[1][0] , \regIn[2][15] , \regIn[2][14] , \regIn[2][13] ,
         \regIn[2][12] , \regIn[2][11] , \regIn[2][10] , \regIn[2][9] ,
         \regIn[2][8] , \regIn[2][7] , \regIn[2][6] , \regIn[2][5] ,
         \regIn[2][4] , \regIn[2][3] , \regIn[2][2] , \regIn[2][1] ,
         \regIn[2][0] , \regIn[3][15] , \regIn[3][14] , \regIn[3][13] ,
         \regIn[3][12] , \regIn[3][11] , \regIn[3][10] , \regIn[3][9] ,
         \regIn[3][8] , \regIn[3][7] , \regIn[3][6] , \regIn[3][5] ,
         \regIn[3][4] , \regIn[3][3] , \regIn[3][2] , \regIn[3][1] ,
         \regIn[3][0] , \regIn[4][15] , \regIn[4][14] , \regIn[4][13] ,
         \regIn[4][12] , \regIn[4][11] , \regIn[4][10] , \regIn[4][9] ,
         \regIn[4][8] , \regIn[4][7] , \regIn[4][6] , \regIn[4][5] ,
         \regIn[4][4] , \regIn[4][3] , \regIn[4][2] , \regIn[4][1] ,
         \regIn[4][0] , \regIn[5][15] , \regIn[5][14] , \regIn[5][13] ,
         \regIn[5][12] , \regIn[5][11] , \regIn[5][10] , \regIn[5][9] ,
         \regIn[5][8] , \regIn[5][7] , \regIn[5][6] , \regIn[5][5] ,
         \regIn[5][4] , \regIn[5][3] , \regIn[5][2] , \regIn[5][1] ,
         \regIn[5][0] , \regIn[6][15] , \regIn[6][14] , \regIn[6][13] ,
         \regIn[6][12] , \regIn[6][11] , \regIn[6][10] , \regIn[6][9] ,
         \regIn[6][8] , \regIn[6][7] , \regIn[6][6] , \regIn[6][5] ,
         \regIn[6][4] , \regIn[6][3] , \regIn[6][2] , \regIn[6][1] ,
         \regIn[6][0] , \regIn[7][15] , \regIn[7][14] , \regIn[7][13] ,
         \regIn[7][12] , \regIn[7][11] , \regIn[7][10] , \regIn[7][9] ,
         \regIn[7][8] , \regIn[7][7] , \regIn[7][6] , \regIn[7][5] ,
         \regIn[7][4] , \regIn[7][3] , \regIn[7][2] , \regIn[7][1] ,
         \regIn[7][0] , \regIn[8][15] , \regIn[8][14] , \regIn[8][13] ,
         \regIn[8][12] , \regIn[8][11] , \regIn[8][10] , \regIn[8][9] ,
         \regIn[8][8] , \regIn[8][7] , \regIn[8][6] , \regIn[8][5] ,
         \regIn[8][4] , \regIn[8][3] , \regIn[8][2] , \regIn[8][1] ,
         \regIn[8][0] , \regIn[9][15] , \regIn[9][14] , \regIn[9][13] ,
         \regIn[9][12] , \regIn[9][11] , \regIn[9][10] , \regIn[9][9] ,
         \regIn[9][8] , \regIn[9][7] , \regIn[9][6] , \regIn[9][5] ,
         \regIn[9][4] , \regIn[9][3] , \regIn[9][2] , \regIn[9][1] ,
         \regIn[9][0] , \regIn[10][15] , \regIn[10][14] , \regIn[10][13] ,
         \regIn[10][12] , \regIn[10][11] , \regIn[10][10] , \regIn[10][9] ,
         \regIn[10][8] , \regIn[10][7] , \regIn[10][6] , \regIn[10][5] ,
         \regIn[10][4] , \regIn[10][3] , \regIn[10][2] , \regIn[10][1] ,
         \regIn[10][0] , \regIn[11][15] , \regIn[11][14] , \regIn[11][13] ,
         \regIn[11][12] , \regIn[11][11] , \regIn[11][10] , \regIn[11][9] ,
         \regIn[11][8] , \regIn[11][7] , \regIn[11][6] , \regIn[11][5] ,
         \regIn[11][4] , \regIn[11][3] , \regIn[11][2] , \regIn[11][1] ,
         \regIn[11][0] , \regIn[12][15] , \regIn[12][14] , \regIn[12][13] ,
         \regIn[12][12] , \regIn[12][11] , \regIn[12][10] , \regIn[12][9] ,
         \regIn[12][8] , \regIn[12][7] , \regIn[12][6] , \regIn[12][5] ,
         \regIn[12][4] , \regIn[12][3] , \regIn[12][2] , \regIn[12][1] ,
         \regIn[12][0] , \regIn[13][15] , \regIn[13][14] , \regIn[13][13] ,
         \regIn[13][12] , \regIn[13][11] , \regIn[13][10] , \regIn[13][9] ,
         \regIn[13][8] , \regIn[13][7] , \regIn[13][6] , \regIn[13][5] ,
         \regIn[13][4] , \regIn[13][3] , \regIn[13][2] , \regIn[13][1] ,
         \regIn[13][0] , \regIn[14][15] , \regIn[14][14] , \regIn[14][13] ,
         \regIn[14][12] , \regIn[14][11] , \regIn[14][10] , \regIn[14][9] ,
         \regIn[14][8] , \regIn[14][7] , \regIn[14][6] , \regIn[14][5] ,
         \regIn[14][4] , \regIn[14][3] , \regIn[14][2] , \regIn[14][1] ,
         \regIn[14][0] , \regIn[15][15] , \regIn[15][14] , \regIn[15][13] ,
         \regIn[15][12] , \regIn[15][11] , \regIn[15][10] , \regIn[15][9] ,
         \regIn[15][8] , \regIn[15][7] , \regIn[15][6] , \regIn[15][5] ,
         \regIn[15][4] , \regIn[15][3] , \regIn[15][2] , \regIn[15][1] ,
         \regIn[15][0] , \regIn[16][15] , \regIn[16][14] , \regIn[16][13] ,
         \regIn[16][12] , \regIn[16][11] , \regIn[16][10] , \regIn[16][9] ,
         \regIn[16][8] , \regIn[16][7] , \regIn[16][6] , \regIn[16][5] ,
         \regIn[16][4] , \regIn[16][3] , \regIn[16][2] , \regIn[16][1] ,
         \regIn[16][0] , \regIn[17][15] , \regIn[17][14] , \regIn[17][13] ,
         \regIn[17][12] , \regIn[17][11] , \regIn[17][10] , \regIn[17][9] ,
         \regIn[17][8] , \regIn[17][7] , \regIn[17][6] , \regIn[17][5] ,
         \regIn[17][4] , \regIn[17][3] , \regIn[17][2] , \regIn[17][1] ,
         \regIn[17][0] , \regIn[18][15] , \regIn[18][14] , \regIn[18][13] ,
         \regIn[18][12] , \regIn[18][11] , \regIn[18][10] , \regIn[18][9] ,
         \regIn[18][8] , \regIn[18][7] , \regIn[18][6] , \regIn[18][5] ,
         \regIn[18][4] , \regIn[18][3] , \regIn[18][2] , \regIn[18][1] ,
         \regIn[18][0] , \regIn[19][15] , \regIn[19][14] , \regIn[19][13] ,
         \regIn[19][12] , \regIn[19][11] , \regIn[19][10] , \regIn[19][9] ,
         \regIn[19][8] , \regIn[19][7] , \regIn[19][6] , \regIn[19][5] ,
         \regIn[19][4] , \regIn[19][3] , \regIn[19][2] , \regIn[19][1] ,
         \regIn[19][0] , \regIn[20][15] , \regIn[20][14] , \regIn[20][13] ,
         \regIn[20][12] , \regIn[20][11] , \regIn[20][10] , \regIn[20][9] ,
         \regIn[20][8] , \regIn[20][7] , \regIn[20][6] , \regIn[20][5] ,
         \regIn[20][4] , \regIn[20][3] , \regIn[20][2] , \regIn[20][1] ,
         \regIn[20][0] , \regIn[21][15] , \regIn[21][14] , \regIn[21][13] ,
         \regIn[21][12] , \regIn[21][11] , \regIn[21][10] , \regIn[21][9] ,
         \regIn[21][8] , \regIn[21][7] , \regIn[21][6] , \regIn[21][5] ,
         \regIn[21][4] , \regIn[21][3] , \regIn[21][2] , \regIn[21][1] ,
         \regIn[21][0] , \regIn[22][15] , \regIn[22][14] , \regIn[22][13] ,
         \regIn[22][12] , \regIn[22][11] , \regIn[22][10] , \regIn[22][9] ,
         \regIn[22][8] , \regIn[22][7] , \regIn[22][6] , \regIn[22][5] ,
         \regIn[22][4] , \regIn[22][3] , \regIn[22][2] , \regIn[22][1] ,
         \regIn[22][0] , \regIn[23][15] , \regIn[23][14] , \regIn[23][13] ,
         \regIn[23][12] , \regIn[23][11] , \regIn[23][10] , \regIn[23][9] ,
         \regIn[23][8] , \regIn[23][7] , \regIn[23][6] , \regIn[23][5] ,
         \regIn[23][4] , \regIn[23][3] , \regIn[23][2] , \regIn[23][1] ,
         \regIn[23][0] , \regIn[24][15] , \regIn[24][14] , \regIn[24][13] ,
         \regIn[24][12] , \regIn[24][11] , \regIn[24][10] , \regIn[24][9] ,
         \regIn[24][8] , \regIn[24][7] , \regIn[24][6] , \regIn[24][5] ,
         \regIn[24][4] , \regIn[24][3] , \regIn[24][2] , \regIn[24][1] ,
         \regIn[24][0] , \regIn[25][15] , \regIn[25][14] , \regIn[25][13] ,
         \regIn[25][12] , \regIn[25][11] , \regIn[25][10] , \regIn[25][9] ,
         \regIn[25][8] , \regIn[25][7] , \regIn[25][6] , \regIn[25][5] ,
         \regIn[25][4] , \regIn[25][3] , \regIn[25][2] , \regIn[25][1] ,
         \regIn[25][0] , \regIn[26][15] , \regIn[26][14] , \regIn[26][13] ,
         \regIn[26][12] , \regIn[26][11] , \regIn[26][10] , \regIn[26][9] ,
         \regIn[26][8] , \regIn[26][7] , \regIn[26][6] , \regIn[26][5] ,
         \regIn[26][4] , \regIn[26][3] , \regIn[26][2] , \regIn[26][1] ,
         \regIn[26][0] , \regIn[27][15] , \regIn[27][14] , \regIn[27][13] ,
         \regIn[27][12] , \regIn[27][11] , \regIn[27][10] , \regIn[27][9] ,
         \regIn[27][8] , \regIn[27][7] , \regIn[27][6] , \regIn[27][5] ,
         \regIn[27][4] , \regIn[27][3] , \regIn[27][2] , \regIn[27][1] ,
         \regIn[27][0] , \regIn[28][15] , \regIn[28][14] , \regIn[28][13] ,
         \regIn[28][12] , \regIn[28][11] , \regIn[28][10] , \regIn[28][9] ,
         \regIn[28][8] , \regIn[28][7] , \regIn[28][6] , \regIn[28][5] ,
         \regIn[28][4] , \regIn[28][3] , \regIn[28][2] , \regIn[28][1] ,
         \regIn[28][0] , \regIn[29][15] , \regIn[29][14] , \regIn[29][13] ,
         \regIn[29][12] , \regIn[29][11] , \regIn[29][10] , \regIn[29][9] ,
         \regIn[29][8] , \regIn[29][7] , \regIn[29][6] , \regIn[29][5] ,
         \regIn[29][4] , \regIn[29][3] , \regIn[29][2] , \regIn[29][1] ,
         \regIn[29][0] , \regIn[30][15] , \regIn[30][14] , \regIn[30][13] ,
         \regIn[30][12] , \regIn[30][11] , \regIn[30][10] , \regIn[30][9] ,
         \regIn[30][8] , \regIn[30][7] , \regIn[30][6] , \regIn[30][5] ,
         \regIn[30][4] , \regIn[30][3] , \regIn[30][2] , \regIn[30][1] ,
         \regIn[30][0] , \regIn[31][15] , \regIn[31][14] , \regIn[31][13] ,
         \regIn[31][12] , \regIn[31][11] , \regIn[31][10] , \regIn[31][9] ,
         \regIn[31][8] , \regIn[31][7] , \regIn[31][6] , \regIn[31][5] ,
         \regIn[31][4] , \regIn[31][3] , \regIn[31][2] , \regIn[31][1] ,
         \regIn[31][0] , N195, N196, N197, N198, N199, N200, N202, N203, N204,
         N205, N206, N207, N208, N209, N210, N211, N212, N213, N215, N216,
         N217, N218, N219, N220, N222, N223, N224, N225, N226, N228, N229,
         N230, N231, N232, N234, N235, N236, N237, N238, N240, N241, N242,
         N243, N244, N245, N247, N248, N249, N250, N251, N253, N254, N255,
         N256, N257, N259, N260, N261, N262, N263, N265, N266, N267, N268,
         N269, N271, N272, N273, N274, N275, N277, N278, N279, N280, N281,
         N283, N284, N285, N286, N287, N289, N290, N291, N292, N293, N296,
         N297, N298, N299, N300, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N314, N315, N316, N317, N318, N320, N321,
         N322, N323, N324, N326, N327, N328, N329, N330, N332, N333, N334,
         N335, N336, N338, N339, N340, N341, N342, N344, N345, N346, N347,
         N348, N350, N351, N352, N353, N354, N356, N357, N358, N359, N360,
         N362, N363, N364, N365, N366, N368, N369, N370, N371, N372, N374,
         N375, N376, N377, N378, N380, N381, N382, N383, N384, N386, N387,
         N388, N389, N390, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69,
         n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83,
         n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97,
         n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109,
         n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120,
         n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142,
         n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153,
         n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164,
         n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175,
         n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186,
         n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197,
         n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208,
         n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219,
         n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230,
         n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241,
         n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252,
         n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263,
         n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285,
         n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
         n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
         n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
         n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802,
         n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813,
         n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824,
         n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835,
         n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
         n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
         n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868,
         n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879,
         n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890,
         n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901,
         n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
         n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923,
         n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934,
         n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945,
         n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956,
         n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967,
         n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978,
         n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
         n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
         n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
         n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020,
         n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030,
         n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040,
         n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050,
         n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060,
         n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070,
         n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080,
         n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090,
         n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100,
         n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110,
         n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120,
         n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130,
         n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140,
         n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150,
         n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160,
         n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
         n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180,
         n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190,
         n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200,
         n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210,
         n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220,
         n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230,
         n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240,
         n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250,
         n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260,
         n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270,
         n1271, n1272, n1273, n1274, n1275;
  assign N208 = addressIn[4];

  INV_X2 I_36 ( .A(N389), .ZN(N390) );
  OR2_X2 C1077 ( .A1(N200), .A2(N388), .ZN(N389) );
  OR2_X2 C1076 ( .A1(N207), .A2(N387), .ZN(N388) );
  OR2_X2 C1075 ( .A1(N220), .A2(N386), .ZN(N387) );
  OR2_X2 C1074 ( .A1(N245), .A2(N307), .ZN(N386) );
  INV_X2 I_35 ( .A(N383), .ZN(N384) );
  OR2_X2 C1065 ( .A1(N207), .A2(N381), .ZN(N382) );
  OR2_X2 C1064 ( .A1(N220), .A2(N380), .ZN(N381) );
  OR2_X2 C1063 ( .A1(N245), .A2(N307), .ZN(N380) );
  INV_X2 I_34 ( .A(N377), .ZN(N378) );
  OR2_X2 C1056 ( .A1(N200), .A2(N376), .ZN(N377) );
  OR2_X2 C1054 ( .A1(N220), .A2(N374), .ZN(N375) );
  OR2_X2 C1053 ( .A1(N245), .A2(N307), .ZN(N374) );
  INV_X2 I_33 ( .A(N371), .ZN(N372) );
  OR2_X2 C1044 ( .A1(N220), .A2(N368), .ZN(N369) );
  OR2_X2 C1043 ( .A1(N245), .A2(N307), .ZN(N368) );
  INV_X2 I_32 ( .A(N365), .ZN(N366) );
  OR2_X2 C1037 ( .A1(N200), .A2(N364), .ZN(N365) );
  OR2_X2 C1036 ( .A1(N207), .A2(N363), .ZN(N364) );
  OR2_X2 C1034 ( .A1(N245), .A2(N307), .ZN(N362) );
  INV_X2 I_31 ( .A(N359), .ZN(N360) );
  OR2_X2 C1026 ( .A1(N207), .A2(N357), .ZN(N358) );
  OR2_X2 C1024 ( .A1(N245), .A2(N307), .ZN(N356) );
  INV_X2 I_30 ( .A(N353), .ZN(N354) );
  OR2_X2 C1018 ( .A1(N200), .A2(N352), .ZN(N353) );
  OR2_X2 C1015 ( .A1(N245), .A2(N307), .ZN(N350) );
  INV_X2 I_29 ( .A(N347), .ZN(N348) );
  OR2_X2 C1006 ( .A1(N245), .A2(N307), .ZN(N344) );
  INV_X2 I_28 ( .A(N341), .ZN(N342) );
  OR2_X2 C1001 ( .A1(N200), .A2(N340), .ZN(N341) );
  OR2_X2 C1000 ( .A1(N207), .A2(N339), .ZN(N340) );
  OR2_X2 C999 ( .A1(N220), .A2(N338), .ZN(N339) );
  INV_X2 I_27 ( .A(N335), .ZN(N336) );
  OR2_X2 C990 ( .A1(N207), .A2(N333), .ZN(N334) );
  OR2_X2 C989 ( .A1(N220), .A2(N332), .ZN(N333) );
  INV_X2 I_26 ( .A(N329), .ZN(N330) );
  OR2_X2 C982 ( .A1(N200), .A2(N328), .ZN(N329) );
  OR2_X2 C980 ( .A1(N220), .A2(N326), .ZN(N327) );
  INV_X2 I_25 ( .A(N323), .ZN(N324) );
  OR2_X2 C971 ( .A1(N220), .A2(N320), .ZN(N321) );
  INV_X2 I_24 ( .A(N317), .ZN(N318) );
  OR2_X2 C965 ( .A1(N200), .A2(N316), .ZN(N317) );
  OR2_X2 C964 ( .A1(N207), .A2(N315), .ZN(N316) );
  INV_X2 I_23 ( .A(N311), .ZN(N312) );
  OR2_X2 C955 ( .A1(N207), .A2(N309), .ZN(N310) );
  INV_X2 I_22 ( .A(N305), .ZN(N306) );
  OR2_X2 C948 ( .A1(N200), .A2(N304), .ZN(N305) );
  INV_X2 I_21 ( .A(N299), .ZN(N300) );
  INV_X2 I_19 ( .A(N292), .ZN(N293) );
  OR2_X2 C933 ( .A1(N200), .A2(N291), .ZN(N292) );
  OR2_X2 C932 ( .A1(N207), .A2(N290), .ZN(N291) );
  OR2_X2 C931 ( .A1(N220), .A2(N289), .ZN(N290) );
  INV_X2 I_18 ( .A(N286), .ZN(N287) );
  OR2_X2 C922 ( .A1(N207), .A2(N284), .ZN(N285) );
  OR2_X2 C921 ( .A1(N220), .A2(N283), .ZN(N284) );
  INV_X2 I_17 ( .A(N280), .ZN(N281) );
  OR2_X2 C914 ( .A1(N200), .A2(N279), .ZN(N280) );
  OR2_X2 C912 ( .A1(N220), .A2(N277), .ZN(N278) );
  INV_X2 I_16 ( .A(N274), .ZN(N275) );
  OR2_X2 C903 ( .A1(N220), .A2(N271), .ZN(N272) );
  INV_X2 I_15 ( .A(N268), .ZN(N269) );
  OR2_X2 C897 ( .A1(N200), .A2(N267), .ZN(N268) );
  OR2_X2 C896 ( .A1(N207), .A2(N266), .ZN(N267) );
  INV_X2 I_14 ( .A(N262), .ZN(N263) );
  OR2_X2 C887 ( .A1(N207), .A2(N260), .ZN(N261) );
  INV_X2 I_13 ( .A(N256), .ZN(N257) );
  OR2_X2 C880 ( .A1(N200), .A2(N255), .ZN(N256) );
  INV_X2 I_12 ( .A(N250), .ZN(N251) );
  INV_X2 I_10 ( .A(N243), .ZN(N244) );
  OR2_X2 C865 ( .A1(N200), .A2(N242), .ZN(N243) );
  OR2_X2 C864 ( .A1(N207), .A2(N241), .ZN(N242) );
  OR2_X2 C863 ( .A1(N220), .A2(N240), .ZN(N241) );
  INV_X2 I_9 ( .A(N237), .ZN(N238) );
  OR2_X2 C855 ( .A1(N207), .A2(N235), .ZN(N236) );
  OR2_X2 C854 ( .A1(N220), .A2(N234), .ZN(N235) );
  INV_X2 I_8 ( .A(N231), .ZN(N232) );
  OR2_X2 C848 ( .A1(N200), .A2(N230), .ZN(N231) );
  OR2_X2 C846 ( .A1(N220), .A2(N228), .ZN(N229) );
  INV_X2 I_7 ( .A(N225), .ZN(N226) );
  OR2_X2 C838 ( .A1(N220), .A2(N222), .ZN(N223) );
  INV_X2 I_5 ( .A(N218), .ZN(N219) );
  OR2_X2 C833 ( .A1(N200), .A2(N217), .ZN(N218) );
  OR2_X2 C832 ( .A1(N207), .A2(N216), .ZN(N217) );
  INV_X2 I_4 ( .A(N212), .ZN(N213) );
  OR2_X2 C824 ( .A1(N207), .A2(N210), .ZN(N211) );
  INV_X2 I_2 ( .A(N205), .ZN(N206) );
  OR2_X2 C818 ( .A1(N200), .A2(N204), .ZN(N205) );
  INV_X2 I_0 ( .A(N198), .ZN(N199) );
  OAI22_X1 U2 ( .A1(n2), .A2(n3), .B1(N257), .B2(n4), .ZN(\regIn[9][9] ) );
  OAI22_X1 U3 ( .A1(n2), .A2(n5), .B1(N257), .B2(n6), .ZN(\regIn[9][8] ) );
  OAI22_X1 U4 ( .A1(n2), .A2(n7), .B1(N257), .B2(n8), .ZN(\regIn[9][7] ) );
  OAI22_X1 U5 ( .A1(n2), .A2(n9), .B1(N257), .B2(n10), .ZN(\regIn[9][6] ) );
  OAI22_X1 U6 ( .A1(n2), .A2(n11), .B1(N257), .B2(n12), .ZN(\regIn[9][5] ) );
  OAI22_X1 U7 ( .A1(n2), .A2(n13), .B1(N257), .B2(n14), .ZN(\regIn[9][4] ) );
  OAI22_X1 U8 ( .A1(n2), .A2(n15), .B1(N257), .B2(n16), .ZN(\regIn[9][3] ) );
  OAI22_X1 U9 ( .A1(n2), .A2(n17), .B1(N257), .B2(n18), .ZN(\regIn[9][2] ) );
  OAI22_X1 U10 ( .A1(n2), .A2(n19), .B1(N257), .B2(n20), .ZN(\regIn[9][1] ) );
  OAI22_X1 U11 ( .A1(n2), .A2(n21), .B1(N257), .B2(n22), .ZN(\regIn[9][15] )
         );
  OAI22_X1 U12 ( .A1(n2), .A2(n23), .B1(N257), .B2(n24), .ZN(\regIn[9][14] )
         );
  OAI22_X1 U13 ( .A1(n2), .A2(n25), .B1(N257), .B2(n26), .ZN(\regIn[9][13] )
         );
  OAI22_X1 U14 ( .A1(n2), .A2(n27), .B1(N257), .B2(n28), .ZN(\regIn[9][12] )
         );
  OAI22_X1 U15 ( .A1(n2), .A2(n29), .B1(N257), .B2(n30), .ZN(\regIn[9][11] )
         );
  OAI22_X1 U16 ( .A1(n2), .A2(n31), .B1(N257), .B2(n32), .ZN(\regIn[9][10] )
         );
  OAI22_X1 U17 ( .A1(n2), .A2(n33), .B1(N257), .B2(n34), .ZN(\regIn[9][0] ) );
  INV_X1 U18 ( .A(N257), .ZN(n2) );
  OAI22_X1 U19 ( .A1(n3), .A2(n35), .B1(N251), .B2(n36), .ZN(\regIn[8][9] ) );
  OAI22_X1 U20 ( .A1(n5), .A2(n35), .B1(N251), .B2(n37), .ZN(\regIn[8][8] ) );
  OAI22_X1 U21 ( .A1(n7), .A2(n35), .B1(N251), .B2(n38), .ZN(\regIn[8][7] ) );
  OAI22_X1 U22 ( .A1(n9), .A2(n35), .B1(N251), .B2(n39), .ZN(\regIn[8][6] ) );
  OAI22_X1 U23 ( .A1(n11), .A2(n35), .B1(N251), .B2(n40), .ZN(\regIn[8][5] )
         );
  OAI22_X1 U24 ( .A1(n13), .A2(n35), .B1(N251), .B2(n41), .ZN(\regIn[8][4] )
         );
  OAI22_X1 U25 ( .A1(n15), .A2(n35), .B1(N251), .B2(n42), .ZN(\regIn[8][3] )
         );
  OAI22_X1 U26 ( .A1(n17), .A2(n35), .B1(N251), .B2(n43), .ZN(\regIn[8][2] )
         );
  OAI22_X1 U27 ( .A1(n19), .A2(n35), .B1(N251), .B2(n44), .ZN(\regIn[8][1] )
         );
  OAI22_X1 U28 ( .A1(n21), .A2(n35), .B1(N251), .B2(n45), .ZN(\regIn[8][15] )
         );
  OAI22_X1 U29 ( .A1(n23), .A2(n35), .B1(N251), .B2(n46), .ZN(\regIn[8][14] )
         );
  OAI22_X1 U30 ( .A1(n25), .A2(n35), .B1(N251), .B2(n47), .ZN(\regIn[8][13] )
         );
  OAI22_X1 U31 ( .A1(n27), .A2(n35), .B1(N251), .B2(n48), .ZN(\regIn[8][12] )
         );
  OAI22_X1 U32 ( .A1(n29), .A2(n35), .B1(N251), .B2(n49), .ZN(\regIn[8][11] )
         );
  OAI22_X1 U33 ( .A1(n31), .A2(n35), .B1(N251), .B2(n50), .ZN(\regIn[8][10] )
         );
  OAI22_X1 U34 ( .A1(n33), .A2(n35), .B1(N251), .B2(n51), .ZN(\regIn[8][0] )
         );
  INV_X1 U35 ( .A(N251), .ZN(n35) );
  INV_X1 U36 ( .A(n52), .ZN(\regIn[7][9] ) );
  AOI22_X1 U37 ( .A1(n1260), .A2(N244), .B1(n53), .B2(\regOut[7][9] ), .ZN(n52) );
  INV_X1 U38 ( .A(n54), .ZN(\regIn[7][8] ) );
  AOI22_X1 U39 ( .A1(n1258), .A2(N244), .B1(n53), .B2(\regOut[7][8] ), .ZN(n54) );
  INV_X1 U40 ( .A(n55), .ZN(\regIn[7][7] ) );
  AOI22_X1 U41 ( .A1(n1256), .A2(N244), .B1(n53), .B2(\regOut[7][7] ), .ZN(n55) );
  INV_X1 U42 ( .A(n56), .ZN(\regIn[7][6] ) );
  AOI22_X1 U43 ( .A1(n1254), .A2(N244), .B1(n53), .B2(\regOut[7][6] ), .ZN(n56) );
  INV_X1 U44 ( .A(n57), .ZN(\regIn[7][5] ) );
  AOI22_X1 U45 ( .A1(n1252), .A2(N244), .B1(n53), .B2(\regOut[7][5] ), .ZN(n57) );
  INV_X1 U46 ( .A(n58), .ZN(\regIn[7][4] ) );
  AOI22_X1 U47 ( .A1(n1253), .A2(N244), .B1(n53), .B2(\regOut[7][4] ), .ZN(n58) );
  INV_X1 U48 ( .A(n59), .ZN(\regIn[7][3] ) );
  AOI22_X1 U49 ( .A1(n1255), .A2(N244), .B1(n53), .B2(\regOut[7][3] ), .ZN(n59) );
  INV_X1 U50 ( .A(n60), .ZN(\regIn[7][2] ) );
  AOI22_X1 U51 ( .A1(n1257), .A2(N244), .B1(n53), .B2(\regOut[7][2] ), .ZN(n60) );
  INV_X1 U52 ( .A(n61), .ZN(\regIn[7][1] ) );
  AOI22_X1 U53 ( .A1(n1259), .A2(N244), .B1(n53), .B2(\regOut[7][1] ), .ZN(n61) );
  INV_X1 U54 ( .A(n62), .ZN(\regIn[7][15] ) );
  AOI22_X1 U55 ( .A1(n1272), .A2(N244), .B1(n53), .B2(\regOut[7][15] ), .ZN(
        n62) );
  INV_X1 U56 ( .A(n63), .ZN(\regIn[7][14] ) );
  AOI22_X1 U57 ( .A1(n1270), .A2(N244), .B1(n53), .B2(\regOut[7][14] ), .ZN(
        n63) );
  INV_X1 U58 ( .A(n64), .ZN(\regIn[7][13] ) );
  AOI22_X1 U59 ( .A1(n1268), .A2(N244), .B1(n53), .B2(\regOut[7][13] ), .ZN(
        n64) );
  INV_X1 U60 ( .A(n65), .ZN(\regIn[7][12] ) );
  AOI22_X1 U61 ( .A1(n1266), .A2(N244), .B1(n53), .B2(\regOut[7][12] ), .ZN(
        n65) );
  INV_X1 U62 ( .A(n66), .ZN(\regIn[7][11] ) );
  AOI22_X1 U63 ( .A1(n1264), .A2(N244), .B1(n53), .B2(\regOut[7][11] ), .ZN(
        n66) );
  INV_X1 U64 ( .A(n67), .ZN(\regIn[7][10] ) );
  AOI22_X1 U65 ( .A1(n1262), .A2(N244), .B1(n53), .B2(\regOut[7][10] ), .ZN(
        n67) );
  INV_X1 U66 ( .A(n68), .ZN(\regIn[7][0] ) );
  AOI22_X1 U67 ( .A1(n1261), .A2(N244), .B1(n53), .B2(\regOut[7][0] ), .ZN(n68) );
  INV_X1 U68 ( .A(N244), .ZN(n53) );
  INV_X1 U69 ( .A(n69), .ZN(\regIn[6][9] ) );
  AOI22_X1 U70 ( .A1(n1260), .A2(N238), .B1(n70), .B2(\regOut[6][9] ), .ZN(n69) );
  INV_X1 U71 ( .A(n71), .ZN(\regIn[6][8] ) );
  AOI22_X1 U72 ( .A1(n1258), .A2(N238), .B1(n70), .B2(\regOut[6][8] ), .ZN(n71) );
  INV_X1 U73 ( .A(n72), .ZN(\regIn[6][7] ) );
  AOI22_X1 U74 ( .A1(n1256), .A2(N238), .B1(n70), .B2(\regOut[6][7] ), .ZN(n72) );
  INV_X1 U75 ( .A(n73), .ZN(\regIn[6][6] ) );
  AOI22_X1 U76 ( .A1(n1254), .A2(N238), .B1(n70), .B2(\regOut[6][6] ), .ZN(n73) );
  INV_X1 U77 ( .A(n74), .ZN(\regIn[6][5] ) );
  AOI22_X1 U78 ( .A1(n1252), .A2(N238), .B1(n70), .B2(\regOut[6][5] ), .ZN(n74) );
  INV_X1 U79 ( .A(n75), .ZN(\regIn[6][4] ) );
  AOI22_X1 U80 ( .A1(n1253), .A2(N238), .B1(n70), .B2(\regOut[6][4] ), .ZN(n75) );
  INV_X1 U81 ( .A(n76), .ZN(\regIn[6][3] ) );
  AOI22_X1 U82 ( .A1(n1255), .A2(N238), .B1(n70), .B2(\regOut[6][3] ), .ZN(n76) );
  INV_X1 U83 ( .A(n77), .ZN(\regIn[6][2] ) );
  AOI22_X1 U84 ( .A1(n1257), .A2(N238), .B1(n70), .B2(\regOut[6][2] ), .ZN(n77) );
  INV_X1 U85 ( .A(n78), .ZN(\regIn[6][1] ) );
  AOI22_X1 U86 ( .A1(n1259), .A2(N238), .B1(n70), .B2(\regOut[6][1] ), .ZN(n78) );
  INV_X1 U87 ( .A(n79), .ZN(\regIn[6][15] ) );
  AOI22_X1 U88 ( .A1(n1272), .A2(N238), .B1(n70), .B2(\regOut[6][15] ), .ZN(
        n79) );
  INV_X1 U89 ( .A(n80), .ZN(\regIn[6][14] ) );
  AOI22_X1 U90 ( .A1(n1270), .A2(N238), .B1(n70), .B2(\regOut[6][14] ), .ZN(
        n80) );
  INV_X1 U91 ( .A(n81), .ZN(\regIn[6][13] ) );
  AOI22_X1 U92 ( .A1(n1268), .A2(N238), .B1(n70), .B2(\regOut[6][13] ), .ZN(
        n81) );
  INV_X1 U93 ( .A(n82), .ZN(\regIn[6][12] ) );
  AOI22_X1 U94 ( .A1(n1266), .A2(N238), .B1(n70), .B2(\regOut[6][12] ), .ZN(
        n82) );
  INV_X1 U95 ( .A(n83), .ZN(\regIn[6][11] ) );
  AOI22_X1 U96 ( .A1(n1264), .A2(N238), .B1(n70), .B2(\regOut[6][11] ), .ZN(
        n83) );
  INV_X1 U97 ( .A(n84), .ZN(\regIn[6][10] ) );
  AOI22_X1 U98 ( .A1(n1262), .A2(N238), .B1(n70), .B2(\regOut[6][10] ), .ZN(
        n84) );
  INV_X1 U99 ( .A(n85), .ZN(\regIn[6][0] ) );
  AOI22_X1 U100 ( .A1(n1261), .A2(N238), .B1(n70), .B2(\regOut[6][0] ), .ZN(
        n85) );
  INV_X1 U101 ( .A(N238), .ZN(n70) );
  OAI22_X1 U102 ( .A1(n3), .A2(n86), .B1(N232), .B2(n87), .ZN(\regIn[5][9] )
         );
  OAI22_X1 U103 ( .A1(n5), .A2(n86), .B1(N232), .B2(n88), .ZN(\regIn[5][8] )
         );
  OAI22_X1 U104 ( .A1(n7), .A2(n86), .B1(N232), .B2(n89), .ZN(\regIn[5][7] )
         );
  OAI22_X1 U105 ( .A1(n9), .A2(n86), .B1(N232), .B2(n90), .ZN(\regIn[5][6] )
         );
  OAI22_X1 U106 ( .A1(n11), .A2(n86), .B1(N232), .B2(n91), .ZN(\regIn[5][5] )
         );
  OAI22_X1 U107 ( .A1(n13), .A2(n86), .B1(N232), .B2(n92), .ZN(\regIn[5][4] )
         );
  OAI22_X1 U108 ( .A1(n15), .A2(n86), .B1(N232), .B2(n93), .ZN(\regIn[5][3] )
         );
  OAI22_X1 U109 ( .A1(n17), .A2(n86), .B1(N232), .B2(n94), .ZN(\regIn[5][2] )
         );
  OAI22_X1 U110 ( .A1(n19), .A2(n86), .B1(N232), .B2(n95), .ZN(\regIn[5][1] )
         );
  OAI22_X1 U111 ( .A1(n21), .A2(n86), .B1(N232), .B2(n96), .ZN(\regIn[5][15] )
         );
  OAI22_X1 U112 ( .A1(n23), .A2(n86), .B1(N232), .B2(n97), .ZN(\regIn[5][14] )
         );
  OAI22_X1 U113 ( .A1(n25), .A2(n86), .B1(N232), .B2(n98), .ZN(\regIn[5][13] )
         );
  OAI22_X1 U114 ( .A1(n27), .A2(n86), .B1(N232), .B2(n99), .ZN(\regIn[5][12] )
         );
  OAI22_X1 U115 ( .A1(n29), .A2(n86), .B1(N232), .B2(n100), .ZN(\regIn[5][11] ) );
  OAI22_X1 U116 ( .A1(n31), .A2(n86), .B1(N232), .B2(n101), .ZN(\regIn[5][10] ) );
  OAI22_X1 U117 ( .A1(n33), .A2(n86), .B1(N232), .B2(n102), .ZN(\regIn[5][0] )
         );
  INV_X1 U118 ( .A(N232), .ZN(n86) );
  OAI22_X1 U119 ( .A1(n3), .A2(n103), .B1(N226), .B2(n104), .ZN(\regIn[4][9] )
         );
  OAI22_X1 U120 ( .A1(n5), .A2(n103), .B1(N226), .B2(n105), .ZN(\regIn[4][8] )
         );
  OAI22_X1 U121 ( .A1(n7), .A2(n103), .B1(N226), .B2(n106), .ZN(\regIn[4][7] )
         );
  OAI22_X1 U122 ( .A1(n9), .A2(n103), .B1(N226), .B2(n107), .ZN(\regIn[4][6] )
         );
  OAI22_X1 U123 ( .A1(n11), .A2(n103), .B1(N226), .B2(n108), .ZN(\regIn[4][5] ) );
  OAI22_X1 U124 ( .A1(n13), .A2(n103), .B1(N226), .B2(n109), .ZN(\regIn[4][4] ) );
  OAI22_X1 U125 ( .A1(n15), .A2(n103), .B1(N226), .B2(n110), .ZN(\regIn[4][3] ) );
  OAI22_X1 U126 ( .A1(n17), .A2(n103), .B1(N226), .B2(n111), .ZN(\regIn[4][2] ) );
  OAI22_X1 U127 ( .A1(n19), .A2(n103), .B1(N226), .B2(n112), .ZN(\regIn[4][1] ) );
  OAI22_X1 U128 ( .A1(n21), .A2(n103), .B1(N226), .B2(n113), .ZN(
        \regIn[4][15] ) );
  OAI22_X1 U129 ( .A1(n23), .A2(n103), .B1(N226), .B2(n114), .ZN(
        \regIn[4][14] ) );
  OAI22_X1 U130 ( .A1(n25), .A2(n103), .B1(N226), .B2(n115), .ZN(
        \regIn[4][13] ) );
  OAI22_X1 U131 ( .A1(n27), .A2(n103), .B1(N226), .B2(n116), .ZN(
        \regIn[4][12] ) );
  OAI22_X1 U132 ( .A1(n29), .A2(n103), .B1(N226), .B2(n117), .ZN(
        \regIn[4][11] ) );
  OAI22_X1 U133 ( .A1(n31), .A2(n103), .B1(N226), .B2(n118), .ZN(
        \regIn[4][10] ) );
  OAI22_X1 U134 ( .A1(n33), .A2(n103), .B1(N226), .B2(n119), .ZN(\regIn[4][0] ) );
  INV_X1 U135 ( .A(N226), .ZN(n103) );
  INV_X1 U136 ( .A(n120), .ZN(\regIn[3][9] ) );
  AOI22_X1 U137 ( .A1(n1260), .A2(N219), .B1(n121), .B2(\regOut[3][9] ), .ZN(
        n120) );
  INV_X1 U138 ( .A(n122), .ZN(\regIn[3][8] ) );
  AOI22_X1 U139 ( .A1(n1258), .A2(N219), .B1(n121), .B2(\regOut[3][8] ), .ZN(
        n122) );
  INV_X1 U140 ( .A(n123), .ZN(\regIn[3][7] ) );
  AOI22_X1 U141 ( .A1(n1256), .A2(N219), .B1(n121), .B2(\regOut[3][7] ), .ZN(
        n123) );
  INV_X1 U142 ( .A(n124), .ZN(\regIn[3][6] ) );
  AOI22_X1 U143 ( .A1(n1254), .A2(N219), .B1(n121), .B2(\regOut[3][6] ), .ZN(
        n124) );
  INV_X1 U144 ( .A(n125), .ZN(\regIn[3][5] ) );
  AOI22_X1 U145 ( .A1(n1252), .A2(N219), .B1(n121), .B2(\regOut[3][5] ), .ZN(
        n125) );
  INV_X1 U146 ( .A(n126), .ZN(\regIn[3][4] ) );
  AOI22_X1 U147 ( .A1(n1253), .A2(N219), .B1(n121), .B2(\regOut[3][4] ), .ZN(
        n126) );
  INV_X1 U148 ( .A(n127), .ZN(\regIn[3][3] ) );
  AOI22_X1 U149 ( .A1(n1255), .A2(N219), .B1(n121), .B2(\regOut[3][3] ), .ZN(
        n127) );
  INV_X1 U150 ( .A(n128), .ZN(\regIn[3][2] ) );
  AOI22_X1 U151 ( .A1(n1257), .A2(N219), .B1(n121), .B2(\regOut[3][2] ), .ZN(
        n128) );
  INV_X1 U152 ( .A(n129), .ZN(\regIn[3][1] ) );
  AOI22_X1 U153 ( .A1(n1259), .A2(N219), .B1(n121), .B2(\regOut[3][1] ), .ZN(
        n129) );
  INV_X1 U154 ( .A(n130), .ZN(\regIn[3][15] ) );
  AOI22_X1 U155 ( .A1(n1272), .A2(N219), .B1(n121), .B2(\regOut[3][15] ), .ZN(
        n130) );
  INV_X1 U156 ( .A(n131), .ZN(\regIn[3][14] ) );
  AOI22_X1 U157 ( .A1(n1270), .A2(N219), .B1(n121), .B2(\regOut[3][14] ), .ZN(
        n131) );
  INV_X1 U158 ( .A(n132), .ZN(\regIn[3][13] ) );
  AOI22_X1 U159 ( .A1(n1268), .A2(N219), .B1(n121), .B2(\regOut[3][13] ), .ZN(
        n132) );
  INV_X1 U160 ( .A(n133), .ZN(\regIn[3][12] ) );
  AOI22_X1 U161 ( .A1(n1266), .A2(N219), .B1(n121), .B2(\regOut[3][12] ), .ZN(
        n133) );
  INV_X1 U162 ( .A(n134), .ZN(\regIn[3][11] ) );
  AOI22_X1 U163 ( .A1(n1264), .A2(N219), .B1(n121), .B2(\regOut[3][11] ), .ZN(
        n134) );
  INV_X1 U164 ( .A(n135), .ZN(\regIn[3][10] ) );
  AOI22_X1 U165 ( .A1(n1262), .A2(N219), .B1(n121), .B2(\regOut[3][10] ), .ZN(
        n135) );
  INV_X1 U166 ( .A(n136), .ZN(\regIn[3][0] ) );
  AOI22_X1 U167 ( .A1(n1261), .A2(N219), .B1(n121), .B2(\regOut[3][0] ), .ZN(
        n136) );
  INV_X1 U168 ( .A(N219), .ZN(n121) );
  OAI22_X1 U169 ( .A1(n3), .A2(n137), .B1(N390), .B2(n138), .ZN(\regIn[31][9] ) );
  OAI22_X1 U170 ( .A1(n5), .A2(n137), .B1(N390), .B2(n139), .ZN(\regIn[31][8] ) );
  OAI22_X1 U171 ( .A1(n7), .A2(n137), .B1(N390), .B2(n140), .ZN(\regIn[31][7] ) );
  OAI22_X1 U172 ( .A1(n9), .A2(n137), .B1(N390), .B2(n141), .ZN(\regIn[31][6] ) );
  OAI22_X1 U173 ( .A1(n11), .A2(n137), .B1(N390), .B2(n142), .ZN(
        \regIn[31][5] ) );
  OAI22_X1 U174 ( .A1(n13), .A2(n137), .B1(N390), .B2(n143), .ZN(
        \regIn[31][4] ) );
  OAI22_X1 U175 ( .A1(n15), .A2(n137), .B1(N390), .B2(n144), .ZN(
        \regIn[31][3] ) );
  OAI22_X1 U176 ( .A1(n17), .A2(n137), .B1(N390), .B2(n145), .ZN(
        \regIn[31][2] ) );
  OAI22_X1 U177 ( .A1(n19), .A2(n137), .B1(N390), .B2(n146), .ZN(
        \regIn[31][1] ) );
  OAI22_X1 U178 ( .A1(n21), .A2(n137), .B1(N390), .B2(n147), .ZN(
        \regIn[31][15] ) );
  OAI22_X1 U179 ( .A1(n23), .A2(n137), .B1(N390), .B2(n148), .ZN(
        \regIn[31][14] ) );
  OAI22_X1 U180 ( .A1(n25), .A2(n137), .B1(N390), .B2(n149), .ZN(
        \regIn[31][13] ) );
  OAI22_X1 U181 ( .A1(n27), .A2(n137), .B1(N390), .B2(n150), .ZN(
        \regIn[31][12] ) );
  OAI22_X1 U182 ( .A1(n29), .A2(n137), .B1(N390), .B2(n151), .ZN(
        \regIn[31][11] ) );
  OAI22_X1 U183 ( .A1(n31), .A2(n137), .B1(N390), .B2(n152), .ZN(
        \regIn[31][10] ) );
  OAI22_X1 U184 ( .A1(n33), .A2(n137), .B1(N390), .B2(n153), .ZN(
        \regIn[31][0] ) );
  INV_X1 U185 ( .A(N390), .ZN(n137) );
  OAI22_X1 U186 ( .A1(n3), .A2(n154), .B1(N384), .B2(n155), .ZN(\regIn[30][9] ) );
  OAI22_X1 U187 ( .A1(n5), .A2(n154), .B1(N384), .B2(n156), .ZN(\regIn[30][8] ) );
  OAI22_X1 U188 ( .A1(n7), .A2(n154), .B1(N384), .B2(n157), .ZN(\regIn[30][7] ) );
  OAI22_X1 U189 ( .A1(n9), .A2(n154), .B1(N384), .B2(n158), .ZN(\regIn[30][6] ) );
  OAI22_X1 U190 ( .A1(n11), .A2(n154), .B1(N384), .B2(n159), .ZN(
        \regIn[30][5] ) );
  OAI22_X1 U191 ( .A1(n13), .A2(n154), .B1(N384), .B2(n160), .ZN(
        \regIn[30][4] ) );
  OAI22_X1 U192 ( .A1(n15), .A2(n154), .B1(N384), .B2(n161), .ZN(
        \regIn[30][3] ) );
  OAI22_X1 U193 ( .A1(n17), .A2(n154), .B1(N384), .B2(n162), .ZN(
        \regIn[30][2] ) );
  OAI22_X1 U194 ( .A1(n19), .A2(n154), .B1(N384), .B2(n163), .ZN(
        \regIn[30][1] ) );
  OAI22_X1 U195 ( .A1(n21), .A2(n154), .B1(N384), .B2(n164), .ZN(
        \regIn[30][15] ) );
  OAI22_X1 U196 ( .A1(n23), .A2(n154), .B1(N384), .B2(n165), .ZN(
        \regIn[30][14] ) );
  OAI22_X1 U197 ( .A1(n25), .A2(n154), .B1(N384), .B2(n166), .ZN(
        \regIn[30][13] ) );
  OAI22_X1 U198 ( .A1(n27), .A2(n154), .B1(N384), .B2(n167), .ZN(
        \regIn[30][12] ) );
  OAI22_X1 U199 ( .A1(n29), .A2(n154), .B1(N384), .B2(n168), .ZN(
        \regIn[30][11] ) );
  OAI22_X1 U200 ( .A1(n31), .A2(n154), .B1(N384), .B2(n169), .ZN(
        \regIn[30][10] ) );
  OAI22_X1 U201 ( .A1(n33), .A2(n154), .B1(N384), .B2(n170), .ZN(
        \regIn[30][0] ) );
  INV_X1 U202 ( .A(N384), .ZN(n154) );
  INV_X1 U203 ( .A(n171), .ZN(\regIn[2][9] ) );
  AOI22_X1 U204 ( .A1(n1260), .A2(N213), .B1(n172), .B2(\regOut[2][9] ), .ZN(
        n171) );
  INV_X1 U205 ( .A(n173), .ZN(\regIn[2][8] ) );
  AOI22_X1 U206 ( .A1(n1258), .A2(N213), .B1(n172), .B2(\regOut[2][8] ), .ZN(
        n173) );
  INV_X1 U207 ( .A(n174), .ZN(\regIn[2][7] ) );
  AOI22_X1 U208 ( .A1(n1256), .A2(N213), .B1(n172), .B2(\regOut[2][7] ), .ZN(
        n174) );
  INV_X1 U209 ( .A(n175), .ZN(\regIn[2][6] ) );
  AOI22_X1 U210 ( .A1(n1254), .A2(N213), .B1(n172), .B2(\regOut[2][6] ), .ZN(
        n175) );
  INV_X1 U211 ( .A(n176), .ZN(\regIn[2][5] ) );
  AOI22_X1 U212 ( .A1(n1252), .A2(N213), .B1(n172), .B2(\regOut[2][5] ), .ZN(
        n176) );
  INV_X1 U213 ( .A(n177), .ZN(\regIn[2][4] ) );
  AOI22_X1 U214 ( .A1(n1253), .A2(N213), .B1(n172), .B2(\regOut[2][4] ), .ZN(
        n177) );
  INV_X1 U215 ( .A(n178), .ZN(\regIn[2][3] ) );
  AOI22_X1 U216 ( .A1(n1255), .A2(N213), .B1(n172), .B2(\regOut[2][3] ), .ZN(
        n178) );
  INV_X1 U217 ( .A(n179), .ZN(\regIn[2][2] ) );
  AOI22_X1 U218 ( .A1(n1257), .A2(N213), .B1(n172), .B2(\regOut[2][2] ), .ZN(
        n179) );
  INV_X1 U219 ( .A(n180), .ZN(\regIn[2][1] ) );
  AOI22_X1 U220 ( .A1(n1259), .A2(N213), .B1(n172), .B2(\regOut[2][1] ), .ZN(
        n180) );
  INV_X1 U221 ( .A(n181), .ZN(\regIn[2][15] ) );
  AOI22_X1 U222 ( .A1(n1272), .A2(N213), .B1(n172), .B2(\regOut[2][15] ), .ZN(
        n181) );
  INV_X1 U223 ( .A(n182), .ZN(\regIn[2][14] ) );
  AOI22_X1 U224 ( .A1(n1270), .A2(N213), .B1(n172), .B2(\regOut[2][14] ), .ZN(
        n182) );
  INV_X1 U225 ( .A(n183), .ZN(\regIn[2][13] ) );
  AOI22_X1 U226 ( .A1(n1268), .A2(N213), .B1(n172), .B2(\regOut[2][13] ), .ZN(
        n183) );
  INV_X1 U227 ( .A(n184), .ZN(\regIn[2][12] ) );
  AOI22_X1 U228 ( .A1(n1266), .A2(N213), .B1(n172), .B2(\regOut[2][12] ), .ZN(
        n184) );
  INV_X1 U229 ( .A(n185), .ZN(\regIn[2][11] ) );
  AOI22_X1 U230 ( .A1(n1264), .A2(N213), .B1(n172), .B2(\regOut[2][11] ), .ZN(
        n185) );
  INV_X1 U231 ( .A(n186), .ZN(\regIn[2][10] ) );
  AOI22_X1 U232 ( .A1(n1262), .A2(N213), .B1(n172), .B2(\regOut[2][10] ), .ZN(
        n186) );
  INV_X1 U233 ( .A(n187), .ZN(\regIn[2][0] ) );
  AOI22_X1 U234 ( .A1(n1261), .A2(N213), .B1(n172), .B2(\regOut[2][0] ), .ZN(
        n187) );
  INV_X1 U235 ( .A(N213), .ZN(n172) );
  INV_X1 U236 ( .A(n188), .ZN(\regIn[29][9] ) );
  AOI22_X1 U237 ( .A1(n1260), .A2(N378), .B1(n189), .B2(\regOut[29][9] ), .ZN(
        n188) );
  INV_X1 U238 ( .A(n190), .ZN(\regIn[29][8] ) );
  AOI22_X1 U239 ( .A1(n1258), .A2(N378), .B1(n189), .B2(\regOut[29][8] ), .ZN(
        n190) );
  INV_X1 U240 ( .A(n191), .ZN(\regIn[29][7] ) );
  AOI22_X1 U241 ( .A1(n1256), .A2(N378), .B1(n189), .B2(\regOut[29][7] ), .ZN(
        n191) );
  INV_X1 U242 ( .A(n192), .ZN(\regIn[29][6] ) );
  AOI22_X1 U243 ( .A1(n1254), .A2(N378), .B1(n189), .B2(\regOut[29][6] ), .ZN(
        n192) );
  INV_X1 U244 ( .A(n193), .ZN(\regIn[29][5] ) );
  AOI22_X1 U245 ( .A1(n1252), .A2(N378), .B1(n189), .B2(\regOut[29][5] ), .ZN(
        n193) );
  INV_X1 U246 ( .A(n194), .ZN(\regIn[29][4] ) );
  AOI22_X1 U247 ( .A1(n1253), .A2(N378), .B1(n189), .B2(\regOut[29][4] ), .ZN(
        n194) );
  INV_X1 U248 ( .A(n195), .ZN(\regIn[29][3] ) );
  AOI22_X1 U249 ( .A1(n1255), .A2(N378), .B1(n189), .B2(\regOut[29][3] ), .ZN(
        n195) );
  INV_X1 U250 ( .A(n196), .ZN(\regIn[29][2] ) );
  AOI22_X1 U251 ( .A1(n1257), .A2(N378), .B1(n189), .B2(\regOut[29][2] ), .ZN(
        n196) );
  INV_X1 U252 ( .A(n197), .ZN(\regIn[29][1] ) );
  AOI22_X1 U253 ( .A1(n1259), .A2(N378), .B1(n189), .B2(\regOut[29][1] ), .ZN(
        n197) );
  INV_X1 U254 ( .A(n198), .ZN(\regIn[29][15] ) );
  AOI22_X1 U255 ( .A1(n1272), .A2(N378), .B1(n189), .B2(\regOut[29][15] ), 
        .ZN(n198) );
  INV_X1 U256 ( .A(n199), .ZN(\regIn[29][14] ) );
  AOI22_X1 U257 ( .A1(n1270), .A2(N378), .B1(n189), .B2(\regOut[29][14] ), 
        .ZN(n199) );
  INV_X1 U258 ( .A(n200), .ZN(\regIn[29][13] ) );
  AOI22_X1 U259 ( .A1(n1268), .A2(N378), .B1(n189), .B2(\regOut[29][13] ), 
        .ZN(n200) );
  INV_X1 U260 ( .A(n201), .ZN(\regIn[29][12] ) );
  AOI22_X1 U261 ( .A1(n1266), .A2(N378), .B1(n189), .B2(\regOut[29][12] ), 
        .ZN(n201) );
  INV_X1 U262 ( .A(n202), .ZN(\regIn[29][11] ) );
  AOI22_X1 U263 ( .A1(n1264), .A2(N378), .B1(n189), .B2(\regOut[29][11] ), 
        .ZN(n202) );
  INV_X1 U264 ( .A(n203), .ZN(\regIn[29][10] ) );
  AOI22_X1 U265 ( .A1(n1262), .A2(N378), .B1(n189), .B2(\regOut[29][10] ), 
        .ZN(n203) );
  INV_X1 U266 ( .A(n204), .ZN(\regIn[29][0] ) );
  AOI22_X1 U267 ( .A1(n1261), .A2(N378), .B1(n189), .B2(\regOut[29][0] ), .ZN(
        n204) );
  INV_X1 U268 ( .A(N378), .ZN(n189) );
  INV_X1 U269 ( .A(n205), .ZN(\regIn[28][9] ) );
  AOI22_X1 U270 ( .A1(n1260), .A2(N372), .B1(n206), .B2(\regOut[28][9] ), .ZN(
        n205) );
  INV_X1 U271 ( .A(n207), .ZN(\regIn[28][8] ) );
  AOI22_X1 U272 ( .A1(n1258), .A2(N372), .B1(n206), .B2(\regOut[28][8] ), .ZN(
        n207) );
  INV_X1 U273 ( .A(n208), .ZN(\regIn[28][7] ) );
  AOI22_X1 U274 ( .A1(n1256), .A2(N372), .B1(n206), .B2(\regOut[28][7] ), .ZN(
        n208) );
  INV_X1 U275 ( .A(n209), .ZN(\regIn[28][6] ) );
  AOI22_X1 U276 ( .A1(n1254), .A2(N372), .B1(n206), .B2(\regOut[28][6] ), .ZN(
        n209) );
  INV_X1 U277 ( .A(n210), .ZN(\regIn[28][5] ) );
  AOI22_X1 U278 ( .A1(n1252), .A2(N372), .B1(n206), .B2(\regOut[28][5] ), .ZN(
        n210) );
  INV_X1 U279 ( .A(n211), .ZN(\regIn[28][4] ) );
  AOI22_X1 U280 ( .A1(n1253), .A2(N372), .B1(n206), .B2(\regOut[28][4] ), .ZN(
        n211) );
  INV_X1 U281 ( .A(n212), .ZN(\regIn[28][3] ) );
  AOI22_X1 U282 ( .A1(n1255), .A2(N372), .B1(n206), .B2(\regOut[28][3] ), .ZN(
        n212) );
  INV_X1 U283 ( .A(n213), .ZN(\regIn[28][2] ) );
  AOI22_X1 U284 ( .A1(n1257), .A2(N372), .B1(n206), .B2(\regOut[28][2] ), .ZN(
        n213) );
  INV_X1 U285 ( .A(n214), .ZN(\regIn[28][1] ) );
  AOI22_X1 U286 ( .A1(n1259), .A2(N372), .B1(n206), .B2(\regOut[28][1] ), .ZN(
        n214) );
  INV_X1 U287 ( .A(n215), .ZN(\regIn[28][15] ) );
  AOI22_X1 U288 ( .A1(n1272), .A2(N372), .B1(n206), .B2(\regOut[28][15] ), 
        .ZN(n215) );
  INV_X1 U289 ( .A(n216), .ZN(\regIn[28][14] ) );
  AOI22_X1 U290 ( .A1(n1270), .A2(N372), .B1(n206), .B2(\regOut[28][14] ), 
        .ZN(n216) );
  INV_X1 U291 ( .A(n217), .ZN(\regIn[28][13] ) );
  AOI22_X1 U292 ( .A1(n1268), .A2(N372), .B1(n206), .B2(\regOut[28][13] ), 
        .ZN(n217) );
  INV_X1 U293 ( .A(n218), .ZN(\regIn[28][12] ) );
  AOI22_X1 U294 ( .A1(n1266), .A2(N372), .B1(n206), .B2(\regOut[28][12] ), 
        .ZN(n218) );
  INV_X1 U295 ( .A(n219), .ZN(\regIn[28][11] ) );
  AOI22_X1 U296 ( .A1(n1264), .A2(N372), .B1(n206), .B2(\regOut[28][11] ), 
        .ZN(n219) );
  INV_X1 U297 ( .A(n220), .ZN(\regIn[28][10] ) );
  AOI22_X1 U298 ( .A1(n1262), .A2(N372), .B1(n206), .B2(\regOut[28][10] ), 
        .ZN(n220) );
  INV_X1 U299 ( .A(n221), .ZN(\regIn[28][0] ) );
  AOI22_X1 U300 ( .A1(n1261), .A2(N372), .B1(n206), .B2(\regOut[28][0] ), .ZN(
        n221) );
  INV_X1 U301 ( .A(N372), .ZN(n206) );
  INV_X1 U302 ( .A(n222), .ZN(\regIn[27][9] ) );
  AOI22_X1 U303 ( .A1(n1260), .A2(N366), .B1(n223), .B2(\regOut[27][9] ), .ZN(
        n222) );
  INV_X1 U304 ( .A(n224), .ZN(\regIn[27][8] ) );
  AOI22_X1 U305 ( .A1(n1258), .A2(N366), .B1(n223), .B2(\regOut[27][8] ), .ZN(
        n224) );
  INV_X1 U306 ( .A(n225), .ZN(\regIn[27][7] ) );
  AOI22_X1 U307 ( .A1(n1256), .A2(N366), .B1(n223), .B2(\regOut[27][7] ), .ZN(
        n225) );
  INV_X1 U308 ( .A(n226), .ZN(\regIn[27][6] ) );
  AOI22_X1 U309 ( .A1(n1254), .A2(N366), .B1(n223), .B2(\regOut[27][6] ), .ZN(
        n226) );
  INV_X1 U310 ( .A(n227), .ZN(\regIn[27][5] ) );
  AOI22_X1 U311 ( .A1(n1252), .A2(N366), .B1(n223), .B2(\regOut[27][5] ), .ZN(
        n227) );
  INV_X1 U312 ( .A(n228), .ZN(\regIn[27][4] ) );
  AOI22_X1 U313 ( .A1(n1253), .A2(N366), .B1(n223), .B2(\regOut[27][4] ), .ZN(
        n228) );
  INV_X1 U314 ( .A(n229), .ZN(\regIn[27][3] ) );
  AOI22_X1 U315 ( .A1(n1255), .A2(N366), .B1(n223), .B2(\regOut[27][3] ), .ZN(
        n229) );
  INV_X1 U316 ( .A(n230), .ZN(\regIn[27][2] ) );
  AOI22_X1 U317 ( .A1(n1257), .A2(N366), .B1(n223), .B2(\regOut[27][2] ), .ZN(
        n230) );
  INV_X1 U318 ( .A(n231), .ZN(\regIn[27][1] ) );
  AOI22_X1 U319 ( .A1(n1259), .A2(N366), .B1(n223), .B2(\regOut[27][1] ), .ZN(
        n231) );
  INV_X1 U320 ( .A(n232), .ZN(\regIn[27][15] ) );
  AOI22_X1 U321 ( .A1(n1272), .A2(N366), .B1(n223), .B2(\regOut[27][15] ), 
        .ZN(n232) );
  INV_X1 U322 ( .A(n233), .ZN(\regIn[27][14] ) );
  AOI22_X1 U323 ( .A1(n1270), .A2(N366), .B1(n223), .B2(\regOut[27][14] ), 
        .ZN(n233) );
  INV_X1 U324 ( .A(n234), .ZN(\regIn[27][13] ) );
  AOI22_X1 U325 ( .A1(n1268), .A2(N366), .B1(n223), .B2(\regOut[27][13] ), 
        .ZN(n234) );
  INV_X1 U326 ( .A(n235), .ZN(\regIn[27][12] ) );
  AOI22_X1 U327 ( .A1(n1266), .A2(N366), .B1(n223), .B2(\regOut[27][12] ), 
        .ZN(n235) );
  INV_X1 U328 ( .A(n236), .ZN(\regIn[27][11] ) );
  AOI22_X1 U329 ( .A1(n1264), .A2(N366), .B1(n223), .B2(\regOut[27][11] ), 
        .ZN(n236) );
  INV_X1 U330 ( .A(n237), .ZN(\regIn[27][10] ) );
  AOI22_X1 U331 ( .A1(n1262), .A2(N366), .B1(n223), .B2(\regOut[27][10] ), 
        .ZN(n237) );
  INV_X1 U332 ( .A(n238), .ZN(\regIn[27][0] ) );
  AOI22_X1 U333 ( .A1(n1261), .A2(N366), .B1(n223), .B2(\regOut[27][0] ), .ZN(
        n238) );
  INV_X1 U334 ( .A(N366), .ZN(n223) );
  INV_X1 U335 ( .A(n239), .ZN(\regIn[26][9] ) );
  AOI22_X1 U336 ( .A1(n1260), .A2(N360), .B1(n240), .B2(\regOut[26][9] ), .ZN(
        n239) );
  INV_X1 U337 ( .A(n241), .ZN(\regIn[26][8] ) );
  AOI22_X1 U338 ( .A1(n1258), .A2(N360), .B1(n240), .B2(\regOut[26][8] ), .ZN(
        n241) );
  INV_X1 U339 ( .A(n242), .ZN(\regIn[26][7] ) );
  AOI22_X1 U340 ( .A1(n1256), .A2(N360), .B1(n240), .B2(\regOut[26][7] ), .ZN(
        n242) );
  INV_X1 U341 ( .A(n243), .ZN(\regIn[26][6] ) );
  AOI22_X1 U342 ( .A1(n1254), .A2(N360), .B1(n240), .B2(\regOut[26][6] ), .ZN(
        n243) );
  INV_X1 U343 ( .A(n244), .ZN(\regIn[26][5] ) );
  AOI22_X1 U344 ( .A1(n1252), .A2(N360), .B1(n240), .B2(\regOut[26][5] ), .ZN(
        n244) );
  INV_X1 U345 ( .A(n245), .ZN(\regIn[26][4] ) );
  AOI22_X1 U346 ( .A1(n1253), .A2(N360), .B1(n240), .B2(\regOut[26][4] ), .ZN(
        n245) );
  INV_X1 U347 ( .A(n246), .ZN(\regIn[26][3] ) );
  AOI22_X1 U348 ( .A1(n1255), .A2(N360), .B1(n240), .B2(\regOut[26][3] ), .ZN(
        n246) );
  INV_X1 U349 ( .A(n247), .ZN(\regIn[26][2] ) );
  AOI22_X1 U350 ( .A1(n1257), .A2(N360), .B1(n240), .B2(\regOut[26][2] ), .ZN(
        n247) );
  INV_X1 U351 ( .A(n248), .ZN(\regIn[26][1] ) );
  AOI22_X1 U352 ( .A1(n1259), .A2(N360), .B1(n240), .B2(\regOut[26][1] ), .ZN(
        n248) );
  INV_X1 U353 ( .A(n249), .ZN(\regIn[26][15] ) );
  AOI22_X1 U354 ( .A1(n1272), .A2(N360), .B1(n240), .B2(\regOut[26][15] ), 
        .ZN(n249) );
  INV_X1 U355 ( .A(n250), .ZN(\regIn[26][14] ) );
  AOI22_X1 U356 ( .A1(n1270), .A2(N360), .B1(n240), .B2(\regOut[26][14] ), 
        .ZN(n250) );
  INV_X1 U357 ( .A(n251), .ZN(\regIn[26][13] ) );
  AOI22_X1 U358 ( .A1(n1268), .A2(N360), .B1(n240), .B2(\regOut[26][13] ), 
        .ZN(n251) );
  INV_X1 U359 ( .A(n252), .ZN(\regIn[26][12] ) );
  AOI22_X1 U360 ( .A1(n1266), .A2(N360), .B1(n240), .B2(\regOut[26][12] ), 
        .ZN(n252) );
  INV_X1 U361 ( .A(n253), .ZN(\regIn[26][11] ) );
  AOI22_X1 U362 ( .A1(n1264), .A2(N360), .B1(n240), .B2(\regOut[26][11] ), 
        .ZN(n253) );
  INV_X1 U363 ( .A(n254), .ZN(\regIn[26][10] ) );
  AOI22_X1 U364 ( .A1(n1262), .A2(N360), .B1(n240), .B2(\regOut[26][10] ), 
        .ZN(n254) );
  INV_X1 U365 ( .A(n255), .ZN(\regIn[26][0] ) );
  AOI22_X1 U366 ( .A1(n1261), .A2(N360), .B1(n240), .B2(\regOut[26][0] ), .ZN(
        n255) );
  INV_X1 U367 ( .A(N360), .ZN(n240) );
  OAI22_X1 U368 ( .A1(n3), .A2(n256), .B1(N354), .B2(n257), .ZN(\regIn[25][9] ) );
  OAI22_X1 U369 ( .A1(n5), .A2(n256), .B1(N354), .B2(n258), .ZN(\regIn[25][8] ) );
  OAI22_X1 U370 ( .A1(n7), .A2(n256), .B1(N354), .B2(n259), .ZN(\regIn[25][7] ) );
  OAI22_X1 U371 ( .A1(n9), .A2(n256), .B1(N354), .B2(n260), .ZN(\regIn[25][6] ) );
  OAI22_X1 U372 ( .A1(n11), .A2(n256), .B1(N354), .B2(n261), .ZN(
        \regIn[25][5] ) );
  OAI22_X1 U373 ( .A1(n13), .A2(n256), .B1(N354), .B2(n262), .ZN(
        \regIn[25][4] ) );
  OAI22_X1 U374 ( .A1(n15), .A2(n256), .B1(N354), .B2(n263), .ZN(
        \regIn[25][3] ) );
  OAI22_X1 U375 ( .A1(n17), .A2(n256), .B1(N354), .B2(n264), .ZN(
        \regIn[25][2] ) );
  OAI22_X1 U376 ( .A1(n19), .A2(n256), .B1(N354), .B2(n265), .ZN(
        \regIn[25][1] ) );
  OAI22_X1 U377 ( .A1(n21), .A2(n256), .B1(N354), .B2(n266), .ZN(
        \regIn[25][15] ) );
  OAI22_X1 U378 ( .A1(n23), .A2(n256), .B1(N354), .B2(n267), .ZN(
        \regIn[25][14] ) );
  OAI22_X1 U379 ( .A1(n25), .A2(n256), .B1(N354), .B2(n268), .ZN(
        \regIn[25][13] ) );
  OAI22_X1 U380 ( .A1(n27), .A2(n256), .B1(N354), .B2(n269), .ZN(
        \regIn[25][12] ) );
  OAI22_X1 U381 ( .A1(n29), .A2(n256), .B1(N354), .B2(n270), .ZN(
        \regIn[25][11] ) );
  OAI22_X1 U382 ( .A1(n31), .A2(n256), .B1(N354), .B2(n271), .ZN(
        \regIn[25][10] ) );
  OAI22_X1 U383 ( .A1(n33), .A2(n256), .B1(N354), .B2(n272), .ZN(
        \regIn[25][0] ) );
  INV_X1 U384 ( .A(N354), .ZN(n256) );
  OAI22_X1 U385 ( .A1(n3), .A2(n273), .B1(N348), .B2(n274), .ZN(\regIn[24][9] ) );
  OAI22_X1 U386 ( .A1(n5), .A2(n273), .B1(N348), .B2(n275), .ZN(\regIn[24][8] ) );
  OAI22_X1 U387 ( .A1(n7), .A2(n273), .B1(N348), .B2(n276), .ZN(\regIn[24][7] ) );
  OAI22_X1 U388 ( .A1(n9), .A2(n273), .B1(N348), .B2(n277), .ZN(\regIn[24][6] ) );
  OAI22_X1 U389 ( .A1(n11), .A2(n273), .B1(N348), .B2(n278), .ZN(
        \regIn[24][5] ) );
  OAI22_X1 U390 ( .A1(n13), .A2(n273), .B1(N348), .B2(n279), .ZN(
        \regIn[24][4] ) );
  OAI22_X1 U391 ( .A1(n15), .A2(n273), .B1(N348), .B2(n280), .ZN(
        \regIn[24][3] ) );
  OAI22_X1 U392 ( .A1(n17), .A2(n273), .B1(N348), .B2(n281), .ZN(
        \regIn[24][2] ) );
  OAI22_X1 U393 ( .A1(n19), .A2(n273), .B1(N348), .B2(n282), .ZN(
        \regIn[24][1] ) );
  OAI22_X1 U394 ( .A1(n21), .A2(n273), .B1(N348), .B2(n283), .ZN(
        \regIn[24][15] ) );
  OAI22_X1 U395 ( .A1(n23), .A2(n273), .B1(N348), .B2(n284), .ZN(
        \regIn[24][14] ) );
  OAI22_X1 U396 ( .A1(n25), .A2(n273), .B1(N348), .B2(n285), .ZN(
        \regIn[24][13] ) );
  OAI22_X1 U397 ( .A1(n27), .A2(n273), .B1(N348), .B2(n286), .ZN(
        \regIn[24][12] ) );
  OAI22_X1 U398 ( .A1(n29), .A2(n273), .B1(N348), .B2(n287), .ZN(
        \regIn[24][11] ) );
  OAI22_X1 U399 ( .A1(n31), .A2(n273), .B1(N348), .B2(n288), .ZN(
        \regIn[24][10] ) );
  OAI22_X1 U400 ( .A1(n33), .A2(n273), .B1(N348), .B2(n289), .ZN(
        \regIn[24][0] ) );
  INV_X1 U401 ( .A(N348), .ZN(n273) );
  INV_X1 U402 ( .A(n290), .ZN(\regIn[23][9] ) );
  AOI22_X1 U403 ( .A1(n1260), .A2(N342), .B1(n291), .B2(\regOut[23][9] ), .ZN(
        n290) );
  INV_X1 U404 ( .A(n292), .ZN(\regIn[23][8] ) );
  AOI22_X1 U405 ( .A1(n1258), .A2(N342), .B1(n291), .B2(\regOut[23][8] ), .ZN(
        n292) );
  INV_X1 U406 ( .A(n293), .ZN(\regIn[23][7] ) );
  AOI22_X1 U407 ( .A1(n1256), .A2(N342), .B1(n291), .B2(\regOut[23][7] ), .ZN(
        n293) );
  INV_X1 U408 ( .A(n294), .ZN(\regIn[23][6] ) );
  AOI22_X1 U409 ( .A1(n1254), .A2(N342), .B1(n291), .B2(\regOut[23][6] ), .ZN(
        n294) );
  INV_X1 U410 ( .A(n295), .ZN(\regIn[23][5] ) );
  AOI22_X1 U411 ( .A1(n1252), .A2(N342), .B1(n291), .B2(\regOut[23][5] ), .ZN(
        n295) );
  INV_X1 U412 ( .A(n296), .ZN(\regIn[23][4] ) );
  AOI22_X1 U413 ( .A1(n1253), .A2(N342), .B1(n291), .B2(\regOut[23][4] ), .ZN(
        n296) );
  INV_X1 U414 ( .A(n297), .ZN(\regIn[23][3] ) );
  AOI22_X1 U415 ( .A1(n1255), .A2(N342), .B1(n291), .B2(\regOut[23][3] ), .ZN(
        n297) );
  INV_X1 U416 ( .A(n298), .ZN(\regIn[23][2] ) );
  AOI22_X1 U417 ( .A1(n1257), .A2(N342), .B1(n291), .B2(\regOut[23][2] ), .ZN(
        n298) );
  INV_X1 U418 ( .A(n299), .ZN(\regIn[23][1] ) );
  AOI22_X1 U419 ( .A1(n1259), .A2(N342), .B1(n291), .B2(\regOut[23][1] ), .ZN(
        n299) );
  INV_X1 U420 ( .A(n300), .ZN(\regIn[23][15] ) );
  AOI22_X1 U421 ( .A1(n1272), .A2(N342), .B1(n291), .B2(\regOut[23][15] ), 
        .ZN(n300) );
  INV_X1 U422 ( .A(n301), .ZN(\regIn[23][14] ) );
  AOI22_X1 U423 ( .A1(n1270), .A2(N342), .B1(n291), .B2(\regOut[23][14] ), 
        .ZN(n301) );
  INV_X1 U424 ( .A(n302), .ZN(\regIn[23][13] ) );
  AOI22_X1 U425 ( .A1(n1268), .A2(N342), .B1(n291), .B2(\regOut[23][13] ), 
        .ZN(n302) );
  INV_X1 U426 ( .A(n303), .ZN(\regIn[23][12] ) );
  AOI22_X1 U427 ( .A1(n1266), .A2(N342), .B1(n291), .B2(\regOut[23][12] ), 
        .ZN(n303) );
  INV_X1 U428 ( .A(n304), .ZN(\regIn[23][11] ) );
  AOI22_X1 U429 ( .A1(n1264), .A2(N342), .B1(n291), .B2(\regOut[23][11] ), 
        .ZN(n304) );
  INV_X1 U430 ( .A(n305), .ZN(\regIn[23][10] ) );
  AOI22_X1 U431 ( .A1(n1262), .A2(N342), .B1(n291), .B2(\regOut[23][10] ), 
        .ZN(n305) );
  INV_X1 U432 ( .A(n306), .ZN(\regIn[23][0] ) );
  AOI22_X1 U433 ( .A1(n1261), .A2(N342), .B1(n291), .B2(\regOut[23][0] ), .ZN(
        n306) );
  INV_X1 U434 ( .A(N342), .ZN(n291) );
  INV_X1 U435 ( .A(n307), .ZN(\regIn[22][9] ) );
  AOI22_X1 U436 ( .A1(n1260), .A2(N336), .B1(n308), .B2(\regOut[22][9] ), .ZN(
        n307) );
  INV_X1 U437 ( .A(n309), .ZN(\regIn[22][8] ) );
  AOI22_X1 U438 ( .A1(n1258), .A2(N336), .B1(n308), .B2(\regOut[22][8] ), .ZN(
        n309) );
  INV_X1 U439 ( .A(n310), .ZN(\regIn[22][7] ) );
  AOI22_X1 U440 ( .A1(n1256), .A2(N336), .B1(n308), .B2(\regOut[22][7] ), .ZN(
        n310) );
  INV_X1 U441 ( .A(n311), .ZN(\regIn[22][6] ) );
  AOI22_X1 U442 ( .A1(n1254), .A2(N336), .B1(n308), .B2(\regOut[22][6] ), .ZN(
        n311) );
  INV_X1 U443 ( .A(n312), .ZN(\regIn[22][5] ) );
  AOI22_X1 U444 ( .A1(n1252), .A2(N336), .B1(n308), .B2(\regOut[22][5] ), .ZN(
        n312) );
  INV_X1 U445 ( .A(n313), .ZN(\regIn[22][4] ) );
  AOI22_X1 U446 ( .A1(n1253), .A2(N336), .B1(n308), .B2(\regOut[22][4] ), .ZN(
        n313) );
  INV_X1 U447 ( .A(n314), .ZN(\regIn[22][3] ) );
  AOI22_X1 U448 ( .A1(n1255), .A2(N336), .B1(n308), .B2(\regOut[22][3] ), .ZN(
        n314) );
  INV_X1 U449 ( .A(n315), .ZN(\regIn[22][2] ) );
  AOI22_X1 U450 ( .A1(n1257), .A2(N336), .B1(n308), .B2(\regOut[22][2] ), .ZN(
        n315) );
  INV_X1 U451 ( .A(n316), .ZN(\regIn[22][1] ) );
  AOI22_X1 U452 ( .A1(n1259), .A2(N336), .B1(n308), .B2(\regOut[22][1] ), .ZN(
        n316) );
  INV_X1 U453 ( .A(n317), .ZN(\regIn[22][15] ) );
  AOI22_X1 U454 ( .A1(n1272), .A2(N336), .B1(n308), .B2(\regOut[22][15] ), 
        .ZN(n317) );
  INV_X1 U455 ( .A(n318), .ZN(\regIn[22][14] ) );
  AOI22_X1 U456 ( .A1(n1270), .A2(N336), .B1(n308), .B2(\regOut[22][14] ), 
        .ZN(n318) );
  INV_X1 U457 ( .A(n319), .ZN(\regIn[22][13] ) );
  AOI22_X1 U458 ( .A1(n1268), .A2(N336), .B1(n308), .B2(\regOut[22][13] ), 
        .ZN(n319) );
  INV_X1 U459 ( .A(n320), .ZN(\regIn[22][12] ) );
  AOI22_X1 U460 ( .A1(n1266), .A2(N336), .B1(n308), .B2(\regOut[22][12] ), 
        .ZN(n320) );
  INV_X1 U461 ( .A(n321), .ZN(\regIn[22][11] ) );
  AOI22_X1 U462 ( .A1(n1264), .A2(N336), .B1(n308), .B2(\regOut[22][11] ), 
        .ZN(n321) );
  INV_X1 U463 ( .A(n322), .ZN(\regIn[22][10] ) );
  AOI22_X1 U464 ( .A1(n1262), .A2(N336), .B1(n308), .B2(\regOut[22][10] ), 
        .ZN(n322) );
  INV_X1 U465 ( .A(n323), .ZN(\regIn[22][0] ) );
  AOI22_X1 U466 ( .A1(n1261), .A2(N336), .B1(n308), .B2(\regOut[22][0] ), .ZN(
        n323) );
  INV_X1 U467 ( .A(N336), .ZN(n308) );
  OAI22_X1 U468 ( .A1(n3), .A2(n324), .B1(N330), .B2(n325), .ZN(\regIn[21][9] ) );
  OAI22_X1 U469 ( .A1(n5), .A2(n324), .B1(N330), .B2(n326), .ZN(\regIn[21][8] ) );
  OAI22_X1 U470 ( .A1(n7), .A2(n324), .B1(N330), .B2(n327), .ZN(\regIn[21][7] ) );
  OAI22_X1 U471 ( .A1(n9), .A2(n324), .B1(N330), .B2(n328), .ZN(\regIn[21][6] ) );
  OAI22_X1 U472 ( .A1(n11), .A2(n324), .B1(N330), .B2(n329), .ZN(
        \regIn[21][5] ) );
  OAI22_X1 U473 ( .A1(n13), .A2(n324), .B1(N330), .B2(n330), .ZN(
        \regIn[21][4] ) );
  OAI22_X1 U474 ( .A1(n15), .A2(n324), .B1(N330), .B2(n331), .ZN(
        \regIn[21][3] ) );
  OAI22_X1 U475 ( .A1(n17), .A2(n324), .B1(N330), .B2(n332), .ZN(
        \regIn[21][2] ) );
  OAI22_X1 U476 ( .A1(n19), .A2(n324), .B1(N330), .B2(n333), .ZN(
        \regIn[21][1] ) );
  OAI22_X1 U477 ( .A1(n21), .A2(n324), .B1(N330), .B2(n334), .ZN(
        \regIn[21][15] ) );
  OAI22_X1 U478 ( .A1(n23), .A2(n324), .B1(N330), .B2(n335), .ZN(
        \regIn[21][14] ) );
  OAI22_X1 U479 ( .A1(n25), .A2(n324), .B1(N330), .B2(n336), .ZN(
        \regIn[21][13] ) );
  OAI22_X1 U480 ( .A1(n27), .A2(n324), .B1(N330), .B2(n337), .ZN(
        \regIn[21][12] ) );
  OAI22_X1 U481 ( .A1(n29), .A2(n324), .B1(N330), .B2(n338), .ZN(
        \regIn[21][11] ) );
  OAI22_X1 U482 ( .A1(n31), .A2(n324), .B1(N330), .B2(n339), .ZN(
        \regIn[21][10] ) );
  OAI22_X1 U483 ( .A1(n33), .A2(n324), .B1(N330), .B2(n340), .ZN(
        \regIn[21][0] ) );
  INV_X1 U484 ( .A(N330), .ZN(n324) );
  OAI22_X1 U485 ( .A1(n3), .A2(n341), .B1(N324), .B2(n342), .ZN(\regIn[20][9] ) );
  OAI22_X1 U486 ( .A1(n5), .A2(n341), .B1(N324), .B2(n343), .ZN(\regIn[20][8] ) );
  OAI22_X1 U487 ( .A1(n7), .A2(n341), .B1(N324), .B2(n344), .ZN(\regIn[20][7] ) );
  OAI22_X1 U488 ( .A1(n9), .A2(n341), .B1(N324), .B2(n345), .ZN(\regIn[20][6] ) );
  OAI22_X1 U489 ( .A1(n11), .A2(n341), .B1(N324), .B2(n346), .ZN(
        \regIn[20][5] ) );
  OAI22_X1 U490 ( .A1(n13), .A2(n341), .B1(N324), .B2(n347), .ZN(
        \regIn[20][4] ) );
  OAI22_X1 U491 ( .A1(n15), .A2(n341), .B1(N324), .B2(n348), .ZN(
        \regIn[20][3] ) );
  OAI22_X1 U492 ( .A1(n17), .A2(n341), .B1(N324), .B2(n349), .ZN(
        \regIn[20][2] ) );
  OAI22_X1 U493 ( .A1(n19), .A2(n341), .B1(N324), .B2(n350), .ZN(
        \regIn[20][1] ) );
  OAI22_X1 U494 ( .A1(n21), .A2(n341), .B1(N324), .B2(n351), .ZN(
        \regIn[20][15] ) );
  OAI22_X1 U495 ( .A1(n23), .A2(n341), .B1(N324), .B2(n352), .ZN(
        \regIn[20][14] ) );
  OAI22_X1 U496 ( .A1(n25), .A2(n341), .B1(N324), .B2(n353), .ZN(
        \regIn[20][13] ) );
  OAI22_X1 U497 ( .A1(n27), .A2(n341), .B1(N324), .B2(n354), .ZN(
        \regIn[20][12] ) );
  OAI22_X1 U498 ( .A1(n29), .A2(n341), .B1(N324), .B2(n355), .ZN(
        \regIn[20][11] ) );
  OAI22_X1 U499 ( .A1(n31), .A2(n341), .B1(N324), .B2(n356), .ZN(
        \regIn[20][10] ) );
  OAI22_X1 U500 ( .A1(n33), .A2(n341), .B1(N324), .B2(n357), .ZN(
        \regIn[20][0] ) );
  INV_X1 U501 ( .A(N324), .ZN(n341) );
  OAI22_X1 U502 ( .A1(n3), .A2(n358), .B1(N206), .B2(n359), .ZN(\regIn[1][9] )
         );
  OAI22_X1 U503 ( .A1(n5), .A2(n358), .B1(N206), .B2(n360), .ZN(\regIn[1][8] )
         );
  OAI22_X1 U504 ( .A1(n7), .A2(n358), .B1(N206), .B2(n361), .ZN(\regIn[1][7] )
         );
  OAI22_X1 U505 ( .A1(n9), .A2(n358), .B1(N206), .B2(n362), .ZN(\regIn[1][6] )
         );
  OAI22_X1 U506 ( .A1(n11), .A2(n358), .B1(N206), .B2(n363), .ZN(\regIn[1][5] ) );
  OAI22_X1 U507 ( .A1(n13), .A2(n358), .B1(N206), .B2(n364), .ZN(\regIn[1][4] ) );
  OAI22_X1 U508 ( .A1(n15), .A2(n358), .B1(N206), .B2(n365), .ZN(\regIn[1][3] ) );
  OAI22_X1 U509 ( .A1(n17), .A2(n358), .B1(N206), .B2(n366), .ZN(\regIn[1][2] ) );
  OAI22_X1 U510 ( .A1(n19), .A2(n358), .B1(N206), .B2(n367), .ZN(\regIn[1][1] ) );
  OAI22_X1 U511 ( .A1(n21), .A2(n358), .B1(N206), .B2(n368), .ZN(
        \regIn[1][15] ) );
  OAI22_X1 U512 ( .A1(n23), .A2(n358), .B1(N206), .B2(n369), .ZN(
        \regIn[1][14] ) );
  OAI22_X1 U513 ( .A1(n25), .A2(n358), .B1(N206), .B2(n370), .ZN(
        \regIn[1][13] ) );
  OAI22_X1 U514 ( .A1(n27), .A2(n358), .B1(N206), .B2(n371), .ZN(
        \regIn[1][12] ) );
  OAI22_X1 U515 ( .A1(n29), .A2(n358), .B1(N206), .B2(n372), .ZN(
        \regIn[1][11] ) );
  OAI22_X1 U516 ( .A1(n31), .A2(n358), .B1(N206), .B2(n373), .ZN(
        \regIn[1][10] ) );
  OAI22_X1 U517 ( .A1(n33), .A2(n358), .B1(N206), .B2(n374), .ZN(\regIn[1][0] ) );
  INV_X1 U518 ( .A(N206), .ZN(n358) );
  INV_X1 U519 ( .A(n375), .ZN(\regIn[19][9] ) );
  AOI22_X1 U520 ( .A1(n1260), .A2(N318), .B1(n376), .B2(\regOut[19][9] ), .ZN(
        n375) );
  INV_X1 U521 ( .A(n377), .ZN(\regIn[19][8] ) );
  AOI22_X1 U522 ( .A1(n1258), .A2(N318), .B1(n376), .B2(\regOut[19][8] ), .ZN(
        n377) );
  INV_X1 U523 ( .A(n378), .ZN(\regIn[19][7] ) );
  AOI22_X1 U524 ( .A1(n1256), .A2(N318), .B1(n376), .B2(\regOut[19][7] ), .ZN(
        n378) );
  INV_X1 U525 ( .A(n379), .ZN(\regIn[19][6] ) );
  AOI22_X1 U526 ( .A1(n1254), .A2(N318), .B1(n376), .B2(\regOut[19][6] ), .ZN(
        n379) );
  INV_X1 U527 ( .A(n380), .ZN(\regIn[19][5] ) );
  AOI22_X1 U528 ( .A1(n1252), .A2(N318), .B1(n376), .B2(\regOut[19][5] ), .ZN(
        n380) );
  INV_X1 U529 ( .A(n381), .ZN(\regIn[19][4] ) );
  AOI22_X1 U530 ( .A1(n1253), .A2(N318), .B1(n376), .B2(\regOut[19][4] ), .ZN(
        n381) );
  INV_X1 U531 ( .A(n382), .ZN(\regIn[19][3] ) );
  AOI22_X1 U532 ( .A1(n1255), .A2(N318), .B1(n376), .B2(\regOut[19][3] ), .ZN(
        n382) );
  INV_X1 U533 ( .A(n383), .ZN(\regIn[19][2] ) );
  AOI22_X1 U534 ( .A1(n1257), .A2(N318), .B1(n376), .B2(\regOut[19][2] ), .ZN(
        n383) );
  INV_X1 U535 ( .A(n384), .ZN(\regIn[19][1] ) );
  AOI22_X1 U536 ( .A1(n1259), .A2(N318), .B1(n376), .B2(\regOut[19][1] ), .ZN(
        n384) );
  INV_X1 U537 ( .A(n385), .ZN(\regIn[19][15] ) );
  AOI22_X1 U538 ( .A1(n1272), .A2(N318), .B1(n376), .B2(\regOut[19][15] ), 
        .ZN(n385) );
  INV_X1 U539 ( .A(n386), .ZN(\regIn[19][14] ) );
  AOI22_X1 U540 ( .A1(n1270), .A2(N318), .B1(n376), .B2(\regOut[19][14] ), 
        .ZN(n386) );
  INV_X1 U541 ( .A(n387), .ZN(\regIn[19][13] ) );
  AOI22_X1 U542 ( .A1(n1268), .A2(N318), .B1(n376), .B2(\regOut[19][13] ), 
        .ZN(n387) );
  INV_X1 U543 ( .A(n388), .ZN(\regIn[19][12] ) );
  AOI22_X1 U544 ( .A1(n1266), .A2(N318), .B1(n376), .B2(\regOut[19][12] ), 
        .ZN(n388) );
  INV_X1 U545 ( .A(n389), .ZN(\regIn[19][11] ) );
  AOI22_X1 U546 ( .A1(n1264), .A2(N318), .B1(n376), .B2(\regOut[19][11] ), 
        .ZN(n389) );
  INV_X1 U547 ( .A(n390), .ZN(\regIn[19][10] ) );
  AOI22_X1 U548 ( .A1(n1262), .A2(N318), .B1(n376), .B2(\regOut[19][10] ), 
        .ZN(n390) );
  INV_X1 U549 ( .A(n391), .ZN(\regIn[19][0] ) );
  AOI22_X1 U550 ( .A1(n1261), .A2(N318), .B1(n376), .B2(\regOut[19][0] ), .ZN(
        n391) );
  INV_X1 U551 ( .A(N318), .ZN(n376) );
  INV_X1 U552 ( .A(n392), .ZN(\regIn[18][9] ) );
  AOI22_X1 U553 ( .A1(n1260), .A2(N312), .B1(n393), .B2(\regOut[18][9] ), .ZN(
        n392) );
  INV_X1 U554 ( .A(n394), .ZN(\regIn[18][8] ) );
  AOI22_X1 U555 ( .A1(n1258), .A2(N312), .B1(n393), .B2(\regOut[18][8] ), .ZN(
        n394) );
  INV_X1 U556 ( .A(n395), .ZN(\regIn[18][7] ) );
  AOI22_X1 U557 ( .A1(n1256), .A2(N312), .B1(n393), .B2(\regOut[18][7] ), .ZN(
        n395) );
  INV_X1 U558 ( .A(n396), .ZN(\regIn[18][6] ) );
  AOI22_X1 U559 ( .A1(n1254), .A2(N312), .B1(n393), .B2(\regOut[18][6] ), .ZN(
        n396) );
  INV_X1 U560 ( .A(n397), .ZN(\regIn[18][5] ) );
  AOI22_X1 U561 ( .A1(n1252), .A2(N312), .B1(n393), .B2(\regOut[18][5] ), .ZN(
        n397) );
  INV_X1 U562 ( .A(n398), .ZN(\regIn[18][4] ) );
  AOI22_X1 U563 ( .A1(n1253), .A2(N312), .B1(n393), .B2(\regOut[18][4] ), .ZN(
        n398) );
  INV_X1 U564 ( .A(n399), .ZN(\regIn[18][3] ) );
  AOI22_X1 U565 ( .A1(n1255), .A2(N312), .B1(n393), .B2(\regOut[18][3] ), .ZN(
        n399) );
  INV_X1 U566 ( .A(n400), .ZN(\regIn[18][2] ) );
  AOI22_X1 U567 ( .A1(n1257), .A2(N312), .B1(n393), .B2(\regOut[18][2] ), .ZN(
        n400) );
  INV_X1 U568 ( .A(n401), .ZN(\regIn[18][1] ) );
  AOI22_X1 U569 ( .A1(n1259), .A2(N312), .B1(n393), .B2(\regOut[18][1] ), .ZN(
        n401) );
  INV_X1 U570 ( .A(n402), .ZN(\regIn[18][15] ) );
  AOI22_X1 U571 ( .A1(n1272), .A2(N312), .B1(n393), .B2(\regOut[18][15] ), 
        .ZN(n402) );
  INV_X1 U572 ( .A(n403), .ZN(\regIn[18][14] ) );
  AOI22_X1 U573 ( .A1(n1270), .A2(N312), .B1(n393), .B2(\regOut[18][14] ), 
        .ZN(n403) );
  INV_X1 U574 ( .A(n404), .ZN(\regIn[18][13] ) );
  AOI22_X1 U575 ( .A1(n1268), .A2(N312), .B1(n393), .B2(\regOut[18][13] ), 
        .ZN(n404) );
  INV_X1 U576 ( .A(n405), .ZN(\regIn[18][12] ) );
  AOI22_X1 U577 ( .A1(n1266), .A2(N312), .B1(n393), .B2(\regOut[18][12] ), 
        .ZN(n405) );
  INV_X1 U578 ( .A(n406), .ZN(\regIn[18][11] ) );
  AOI22_X1 U579 ( .A1(n1264), .A2(N312), .B1(n393), .B2(\regOut[18][11] ), 
        .ZN(n406) );
  INV_X1 U580 ( .A(n407), .ZN(\regIn[18][10] ) );
  AOI22_X1 U581 ( .A1(n1262), .A2(N312), .B1(n393), .B2(\regOut[18][10] ), 
        .ZN(n407) );
  INV_X1 U582 ( .A(n408), .ZN(\regIn[18][0] ) );
  AOI22_X1 U583 ( .A1(n1261), .A2(N312), .B1(n393), .B2(\regOut[18][0] ), .ZN(
        n408) );
  INV_X1 U584 ( .A(N312), .ZN(n393) );
  OAI22_X1 U585 ( .A1(n3), .A2(n409), .B1(N306), .B2(n410), .ZN(\regIn[17][9] ) );
  OAI22_X1 U586 ( .A1(n5), .A2(n409), .B1(N306), .B2(n411), .ZN(\regIn[17][8] ) );
  OAI22_X1 U587 ( .A1(n7), .A2(n409), .B1(N306), .B2(n412), .ZN(\regIn[17][7] ) );
  OAI22_X1 U588 ( .A1(n9), .A2(n409), .B1(N306), .B2(n413), .ZN(\regIn[17][6] ) );
  OAI22_X1 U589 ( .A1(n11), .A2(n409), .B1(N306), .B2(n414), .ZN(
        \regIn[17][5] ) );
  OAI22_X1 U590 ( .A1(n13), .A2(n409), .B1(N306), .B2(n415), .ZN(
        \regIn[17][4] ) );
  OAI22_X1 U591 ( .A1(n15), .A2(n409), .B1(N306), .B2(n416), .ZN(
        \regIn[17][3] ) );
  OAI22_X1 U592 ( .A1(n17), .A2(n409), .B1(N306), .B2(n417), .ZN(
        \regIn[17][2] ) );
  OAI22_X1 U593 ( .A1(n19), .A2(n409), .B1(N306), .B2(n418), .ZN(
        \regIn[17][1] ) );
  OAI22_X1 U594 ( .A1(n21), .A2(n409), .B1(N306), .B2(n419), .ZN(
        \regIn[17][15] ) );
  OAI22_X1 U595 ( .A1(n23), .A2(n409), .B1(N306), .B2(n420), .ZN(
        \regIn[17][14] ) );
  OAI22_X1 U596 ( .A1(n25), .A2(n409), .B1(N306), .B2(n421), .ZN(
        \regIn[17][13] ) );
  OAI22_X1 U597 ( .A1(n27), .A2(n409), .B1(N306), .B2(n422), .ZN(
        \regIn[17][12] ) );
  OAI22_X1 U598 ( .A1(n29), .A2(n409), .B1(N306), .B2(n423), .ZN(
        \regIn[17][11] ) );
  OAI22_X1 U599 ( .A1(n31), .A2(n409), .B1(N306), .B2(n424), .ZN(
        \regIn[17][10] ) );
  OAI22_X1 U600 ( .A1(n33), .A2(n409), .B1(N306), .B2(n425), .ZN(
        \regIn[17][0] ) );
  INV_X1 U601 ( .A(N306), .ZN(n409) );
  OAI22_X1 U602 ( .A1(n3), .A2(n426), .B1(N300), .B2(n427), .ZN(\regIn[16][9] ) );
  OAI22_X1 U603 ( .A1(n5), .A2(n426), .B1(N300), .B2(n428), .ZN(\regIn[16][8] ) );
  OAI22_X1 U604 ( .A1(n7), .A2(n426), .B1(N300), .B2(n429), .ZN(\regIn[16][7] ) );
  OAI22_X1 U605 ( .A1(n9), .A2(n426), .B1(N300), .B2(n430), .ZN(\regIn[16][6] ) );
  OAI22_X1 U606 ( .A1(n11), .A2(n426), .B1(N300), .B2(n431), .ZN(
        \regIn[16][5] ) );
  OAI22_X1 U607 ( .A1(n13), .A2(n426), .B1(N300), .B2(n432), .ZN(
        \regIn[16][4] ) );
  OAI22_X1 U608 ( .A1(n15), .A2(n426), .B1(N300), .B2(n433), .ZN(
        \regIn[16][3] ) );
  OAI22_X1 U609 ( .A1(n17), .A2(n426), .B1(N300), .B2(n434), .ZN(
        \regIn[16][2] ) );
  OAI22_X1 U610 ( .A1(n19), .A2(n426), .B1(N300), .B2(n435), .ZN(
        \regIn[16][1] ) );
  OAI22_X1 U611 ( .A1(n21), .A2(n426), .B1(N300), .B2(n436), .ZN(
        \regIn[16][15] ) );
  OAI22_X1 U612 ( .A1(n23), .A2(n426), .B1(N300), .B2(n437), .ZN(
        \regIn[16][14] ) );
  OAI22_X1 U613 ( .A1(n25), .A2(n426), .B1(N300), .B2(n438), .ZN(
        \regIn[16][13] ) );
  OAI22_X1 U614 ( .A1(n27), .A2(n426), .B1(N300), .B2(n439), .ZN(
        \regIn[16][12] ) );
  OAI22_X1 U615 ( .A1(n29), .A2(n426), .B1(N300), .B2(n440), .ZN(
        \regIn[16][11] ) );
  OAI22_X1 U616 ( .A1(n31), .A2(n426), .B1(N300), .B2(n441), .ZN(
        \regIn[16][10] ) );
  OAI22_X1 U617 ( .A1(n33), .A2(n426), .B1(N300), .B2(n442), .ZN(
        \regIn[16][0] ) );
  INV_X1 U618 ( .A(N300), .ZN(n426) );
  INV_X1 U619 ( .A(n443), .ZN(\regIn[15][9] ) );
  AOI22_X1 U620 ( .A1(n1260), .A2(N293), .B1(n444), .B2(\regOut[15][9] ), .ZN(
        n443) );
  INV_X1 U621 ( .A(n445), .ZN(\regIn[15][8] ) );
  AOI22_X1 U622 ( .A1(n1258), .A2(N293), .B1(n444), .B2(\regOut[15][8] ), .ZN(
        n445) );
  INV_X1 U623 ( .A(n446), .ZN(\regIn[15][7] ) );
  AOI22_X1 U624 ( .A1(n1256), .A2(N293), .B1(n444), .B2(\regOut[15][7] ), .ZN(
        n446) );
  INV_X1 U625 ( .A(n447), .ZN(\regIn[15][6] ) );
  AOI22_X1 U626 ( .A1(n1254), .A2(N293), .B1(n444), .B2(\regOut[15][6] ), .ZN(
        n447) );
  INV_X1 U627 ( .A(n448), .ZN(\regIn[15][5] ) );
  AOI22_X1 U628 ( .A1(n1252), .A2(N293), .B1(n444), .B2(\regOut[15][5] ), .ZN(
        n448) );
  INV_X1 U629 ( .A(n449), .ZN(\regIn[15][4] ) );
  AOI22_X1 U630 ( .A1(n1253), .A2(N293), .B1(n444), .B2(\regOut[15][4] ), .ZN(
        n449) );
  INV_X1 U631 ( .A(n450), .ZN(\regIn[15][3] ) );
  AOI22_X1 U632 ( .A1(n1255), .A2(N293), .B1(n444), .B2(\regOut[15][3] ), .ZN(
        n450) );
  INV_X1 U633 ( .A(n451), .ZN(\regIn[15][2] ) );
  AOI22_X1 U634 ( .A1(n1257), .A2(N293), .B1(n444), .B2(\regOut[15][2] ), .ZN(
        n451) );
  INV_X1 U635 ( .A(n452), .ZN(\regIn[15][1] ) );
  AOI22_X1 U636 ( .A1(n1259), .A2(N293), .B1(n444), .B2(\regOut[15][1] ), .ZN(
        n452) );
  INV_X1 U637 ( .A(n453), .ZN(\regIn[15][15] ) );
  AOI22_X1 U638 ( .A1(n1272), .A2(N293), .B1(n444), .B2(\regOut[15][15] ), 
        .ZN(n453) );
  INV_X1 U639 ( .A(n454), .ZN(\regIn[15][14] ) );
  AOI22_X1 U640 ( .A1(n1270), .A2(N293), .B1(n444), .B2(\regOut[15][14] ), 
        .ZN(n454) );
  INV_X1 U641 ( .A(n455), .ZN(\regIn[15][13] ) );
  AOI22_X1 U642 ( .A1(n1268), .A2(N293), .B1(n444), .B2(\regOut[15][13] ), 
        .ZN(n455) );
  INV_X1 U643 ( .A(n456), .ZN(\regIn[15][12] ) );
  AOI22_X1 U644 ( .A1(n1266), .A2(N293), .B1(n444), .B2(\regOut[15][12] ), 
        .ZN(n456) );
  INV_X1 U645 ( .A(n457), .ZN(\regIn[15][11] ) );
  AOI22_X1 U646 ( .A1(n1264), .A2(N293), .B1(n444), .B2(\regOut[15][11] ), 
        .ZN(n457) );
  INV_X1 U647 ( .A(n458), .ZN(\regIn[15][10] ) );
  AOI22_X1 U648 ( .A1(n1262), .A2(N293), .B1(n444), .B2(\regOut[15][10] ), 
        .ZN(n458) );
  INV_X1 U649 ( .A(n459), .ZN(\regIn[15][0] ) );
  AOI22_X1 U650 ( .A1(n1261), .A2(N293), .B1(n444), .B2(\regOut[15][0] ), .ZN(
        n459) );
  INV_X1 U651 ( .A(N293), .ZN(n444) );
  INV_X1 U652 ( .A(n460), .ZN(\regIn[14][9] ) );
  AOI22_X1 U653 ( .A1(n1260), .A2(N287), .B1(n461), .B2(\regOut[14][9] ), .ZN(
        n460) );
  INV_X1 U654 ( .A(n462), .ZN(\regIn[14][8] ) );
  AOI22_X1 U655 ( .A1(n1258), .A2(N287), .B1(n461), .B2(\regOut[14][8] ), .ZN(
        n462) );
  INV_X1 U656 ( .A(n463), .ZN(\regIn[14][7] ) );
  AOI22_X1 U657 ( .A1(n1256), .A2(N287), .B1(n461), .B2(\regOut[14][7] ), .ZN(
        n463) );
  INV_X1 U658 ( .A(n464), .ZN(\regIn[14][6] ) );
  AOI22_X1 U659 ( .A1(n1254), .A2(N287), .B1(n461), .B2(\regOut[14][6] ), .ZN(
        n464) );
  INV_X1 U660 ( .A(n465), .ZN(\regIn[14][5] ) );
  AOI22_X1 U661 ( .A1(n1252), .A2(N287), .B1(n461), .B2(\regOut[14][5] ), .ZN(
        n465) );
  INV_X1 U662 ( .A(n466), .ZN(\regIn[14][4] ) );
  AOI22_X1 U663 ( .A1(n1253), .A2(N287), .B1(n461), .B2(\regOut[14][4] ), .ZN(
        n466) );
  INV_X1 U664 ( .A(n467), .ZN(\regIn[14][3] ) );
  AOI22_X1 U665 ( .A1(n1255), .A2(N287), .B1(n461), .B2(\regOut[14][3] ), .ZN(
        n467) );
  INV_X1 U666 ( .A(n468), .ZN(\regIn[14][2] ) );
  AOI22_X1 U667 ( .A1(n1257), .A2(N287), .B1(n461), .B2(\regOut[14][2] ), .ZN(
        n468) );
  INV_X1 U668 ( .A(n469), .ZN(\regIn[14][1] ) );
  AOI22_X1 U669 ( .A1(n1259), .A2(N287), .B1(n461), .B2(\regOut[14][1] ), .ZN(
        n469) );
  INV_X1 U670 ( .A(n470), .ZN(\regIn[14][15] ) );
  AOI22_X1 U671 ( .A1(n1272), .A2(N287), .B1(n461), .B2(\regOut[14][15] ), 
        .ZN(n470) );
  INV_X1 U672 ( .A(n471), .ZN(\regIn[14][14] ) );
  AOI22_X1 U673 ( .A1(n1270), .A2(N287), .B1(n461), .B2(\regOut[14][14] ), 
        .ZN(n471) );
  INV_X1 U674 ( .A(n472), .ZN(\regIn[14][13] ) );
  AOI22_X1 U675 ( .A1(n1268), .A2(N287), .B1(n461), .B2(\regOut[14][13] ), 
        .ZN(n472) );
  INV_X1 U676 ( .A(n473), .ZN(\regIn[14][12] ) );
  AOI22_X1 U677 ( .A1(n1266), .A2(N287), .B1(n461), .B2(\regOut[14][12] ), 
        .ZN(n473) );
  INV_X1 U678 ( .A(n474), .ZN(\regIn[14][11] ) );
  AOI22_X1 U679 ( .A1(n1264), .A2(N287), .B1(n461), .B2(\regOut[14][11] ), 
        .ZN(n474) );
  INV_X1 U680 ( .A(n475), .ZN(\regIn[14][10] ) );
  AOI22_X1 U681 ( .A1(n1262), .A2(N287), .B1(n461), .B2(\regOut[14][10] ), 
        .ZN(n475) );
  INV_X1 U682 ( .A(n476), .ZN(\regIn[14][0] ) );
  AOI22_X1 U683 ( .A1(n1261), .A2(N287), .B1(n461), .B2(\regOut[14][0] ), .ZN(
        n476) );
  INV_X1 U684 ( .A(N287), .ZN(n461) );
  OAI22_X1 U685 ( .A1(n3), .A2(n477), .B1(N281), .B2(n478), .ZN(\regIn[13][9] ) );
  OAI22_X1 U686 ( .A1(n5), .A2(n477), .B1(N281), .B2(n479), .ZN(\regIn[13][8] ) );
  OAI22_X1 U687 ( .A1(n7), .A2(n477), .B1(N281), .B2(n480), .ZN(\regIn[13][7] ) );
  OAI22_X1 U688 ( .A1(n9), .A2(n477), .B1(N281), .B2(n481), .ZN(\regIn[13][6] ) );
  OAI22_X1 U689 ( .A1(n11), .A2(n477), .B1(N281), .B2(n482), .ZN(
        \regIn[13][5] ) );
  OAI22_X1 U690 ( .A1(n13), .A2(n477), .B1(N281), .B2(n483), .ZN(
        \regIn[13][4] ) );
  OAI22_X1 U691 ( .A1(n15), .A2(n477), .B1(N281), .B2(n484), .ZN(
        \regIn[13][3] ) );
  OAI22_X1 U692 ( .A1(n17), .A2(n477), .B1(N281), .B2(n485), .ZN(
        \regIn[13][2] ) );
  OAI22_X1 U693 ( .A1(n19), .A2(n477), .B1(N281), .B2(n486), .ZN(
        \regIn[13][1] ) );
  OAI22_X1 U694 ( .A1(n21), .A2(n477), .B1(N281), .B2(n487), .ZN(
        \regIn[13][15] ) );
  OAI22_X1 U695 ( .A1(n23), .A2(n477), .B1(N281), .B2(n488), .ZN(
        \regIn[13][14] ) );
  OAI22_X1 U696 ( .A1(n25), .A2(n477), .B1(N281), .B2(n489), .ZN(
        \regIn[13][13] ) );
  OAI22_X1 U697 ( .A1(n27), .A2(n477), .B1(N281), .B2(n490), .ZN(
        \regIn[13][12] ) );
  OAI22_X1 U698 ( .A1(n29), .A2(n477), .B1(N281), .B2(n491), .ZN(
        \regIn[13][11] ) );
  OAI22_X1 U699 ( .A1(n31), .A2(n477), .B1(N281), .B2(n492), .ZN(
        \regIn[13][10] ) );
  OAI22_X1 U700 ( .A1(n33), .A2(n477), .B1(N281), .B2(n493), .ZN(
        \regIn[13][0] ) );
  INV_X1 U701 ( .A(N281), .ZN(n477) );
  OAI22_X1 U702 ( .A1(n3), .A2(n494), .B1(N275), .B2(n495), .ZN(\regIn[12][9] ) );
  OAI22_X1 U703 ( .A1(n5), .A2(n494), .B1(N275), .B2(n496), .ZN(\regIn[12][8] ) );
  OAI22_X1 U704 ( .A1(n7), .A2(n494), .B1(N275), .B2(n497), .ZN(\regIn[12][7] ) );
  OAI22_X1 U705 ( .A1(n9), .A2(n494), .B1(N275), .B2(n498), .ZN(\regIn[12][6] ) );
  OAI22_X1 U706 ( .A1(n11), .A2(n494), .B1(N275), .B2(n499), .ZN(
        \regIn[12][5] ) );
  OAI22_X1 U707 ( .A1(n13), .A2(n494), .B1(N275), .B2(n500), .ZN(
        \regIn[12][4] ) );
  OAI22_X1 U708 ( .A1(n15), .A2(n494), .B1(N275), .B2(n501), .ZN(
        \regIn[12][3] ) );
  OAI22_X1 U709 ( .A1(n17), .A2(n494), .B1(N275), .B2(n502), .ZN(
        \regIn[12][2] ) );
  OAI22_X1 U710 ( .A1(n19), .A2(n494), .B1(N275), .B2(n503), .ZN(
        \regIn[12][1] ) );
  OAI22_X1 U711 ( .A1(n21), .A2(n494), .B1(N275), .B2(n504), .ZN(
        \regIn[12][15] ) );
  OAI22_X1 U712 ( .A1(n23), .A2(n494), .B1(N275), .B2(n505), .ZN(
        \regIn[12][14] ) );
  OAI22_X1 U713 ( .A1(n25), .A2(n494), .B1(N275), .B2(n506), .ZN(
        \regIn[12][13] ) );
  OAI22_X1 U714 ( .A1(n27), .A2(n494), .B1(N275), .B2(n507), .ZN(
        \regIn[12][12] ) );
  OAI22_X1 U715 ( .A1(n29), .A2(n494), .B1(N275), .B2(n508), .ZN(
        \regIn[12][11] ) );
  OAI22_X1 U716 ( .A1(n31), .A2(n494), .B1(N275), .B2(n509), .ZN(
        \regIn[12][10] ) );
  OAI22_X1 U717 ( .A1(n33), .A2(n494), .B1(N275), .B2(n510), .ZN(
        \regIn[12][0] ) );
  INV_X1 U718 ( .A(N275), .ZN(n494) );
  INV_X1 U719 ( .A(n511), .ZN(\regIn[11][9] ) );
  AOI22_X1 U720 ( .A1(n1260), .A2(N269), .B1(n512), .B2(\regOut[11][9] ), .ZN(
        n511) );
  INV_X1 U721 ( .A(n513), .ZN(\regIn[11][8] ) );
  AOI22_X1 U722 ( .A1(n1258), .A2(N269), .B1(n512), .B2(\regOut[11][8] ), .ZN(
        n513) );
  INV_X1 U723 ( .A(n514), .ZN(\regIn[11][7] ) );
  AOI22_X1 U724 ( .A1(n1256), .A2(N269), .B1(n512), .B2(\regOut[11][7] ), .ZN(
        n514) );
  INV_X1 U725 ( .A(n515), .ZN(\regIn[11][6] ) );
  AOI22_X1 U726 ( .A1(n1254), .A2(N269), .B1(n512), .B2(\regOut[11][6] ), .ZN(
        n515) );
  INV_X1 U727 ( .A(n516), .ZN(\regIn[11][5] ) );
  AOI22_X1 U728 ( .A1(n1252), .A2(N269), .B1(n512), .B2(\regOut[11][5] ), .ZN(
        n516) );
  INV_X1 U729 ( .A(n517), .ZN(\regIn[11][4] ) );
  AOI22_X1 U730 ( .A1(n1253), .A2(N269), .B1(n512), .B2(\regOut[11][4] ), .ZN(
        n517) );
  INV_X1 U731 ( .A(n518), .ZN(\regIn[11][3] ) );
  AOI22_X1 U732 ( .A1(n1255), .A2(N269), .B1(n512), .B2(\regOut[11][3] ), .ZN(
        n518) );
  INV_X1 U733 ( .A(n519), .ZN(\regIn[11][2] ) );
  AOI22_X1 U734 ( .A1(n1257), .A2(N269), .B1(n512), .B2(\regOut[11][2] ), .ZN(
        n519) );
  INV_X1 U735 ( .A(n520), .ZN(\regIn[11][1] ) );
  AOI22_X1 U736 ( .A1(n1259), .A2(N269), .B1(n512), .B2(\regOut[11][1] ), .ZN(
        n520) );
  INV_X1 U737 ( .A(n521), .ZN(\regIn[11][15] ) );
  AOI22_X1 U738 ( .A1(n1272), .A2(N269), .B1(n512), .B2(\regOut[11][15] ), 
        .ZN(n521) );
  INV_X1 U739 ( .A(n522), .ZN(\regIn[11][14] ) );
  AOI22_X1 U740 ( .A1(n1270), .A2(N269), .B1(n512), .B2(\regOut[11][14] ), 
        .ZN(n522) );
  INV_X1 U741 ( .A(n523), .ZN(\regIn[11][13] ) );
  AOI22_X1 U742 ( .A1(n1268), .A2(N269), .B1(n512), .B2(\regOut[11][13] ), 
        .ZN(n523) );
  INV_X1 U743 ( .A(n524), .ZN(\regIn[11][12] ) );
  AOI22_X1 U744 ( .A1(n1266), .A2(N269), .B1(n512), .B2(\regOut[11][12] ), 
        .ZN(n524) );
  INV_X1 U745 ( .A(n525), .ZN(\regIn[11][11] ) );
  AOI22_X1 U746 ( .A1(n1264), .A2(N269), .B1(n512), .B2(\regOut[11][11] ), 
        .ZN(n525) );
  INV_X1 U747 ( .A(n526), .ZN(\regIn[11][10] ) );
  AOI22_X1 U748 ( .A1(n1262), .A2(N269), .B1(n512), .B2(\regOut[11][10] ), 
        .ZN(n526) );
  INV_X1 U749 ( .A(n527), .ZN(\regIn[11][0] ) );
  AOI22_X1 U750 ( .A1(n1261), .A2(N269), .B1(n512), .B2(\regOut[11][0] ), .ZN(
        n527) );
  INV_X1 U751 ( .A(N269), .ZN(n512) );
  INV_X1 U752 ( .A(n528), .ZN(\regIn[10][9] ) );
  AOI22_X1 U753 ( .A1(n1260), .A2(N263), .B1(n529), .B2(\regOut[10][9] ), .ZN(
        n528) );
  INV_X1 U754 ( .A(n530), .ZN(\regIn[10][8] ) );
  AOI22_X1 U755 ( .A1(n1258), .A2(N263), .B1(n529), .B2(\regOut[10][8] ), .ZN(
        n530) );
  INV_X1 U756 ( .A(n531), .ZN(\regIn[10][7] ) );
  AOI22_X1 U757 ( .A1(n1256), .A2(N263), .B1(n529), .B2(\regOut[10][7] ), .ZN(
        n531) );
  INV_X1 U758 ( .A(n532), .ZN(\regIn[10][6] ) );
  AOI22_X1 U759 ( .A1(n1254), .A2(N263), .B1(n529), .B2(\regOut[10][6] ), .ZN(
        n532) );
  INV_X1 U760 ( .A(n533), .ZN(\regIn[10][5] ) );
  AOI22_X1 U761 ( .A1(n1252), .A2(N263), .B1(n529), .B2(\regOut[10][5] ), .ZN(
        n533) );
  INV_X1 U762 ( .A(n534), .ZN(\regIn[10][4] ) );
  AOI22_X1 U763 ( .A1(n1253), .A2(N263), .B1(n529), .B2(\regOut[10][4] ), .ZN(
        n534) );
  INV_X1 U764 ( .A(n535), .ZN(\regIn[10][3] ) );
  AOI22_X1 U765 ( .A1(n1255), .A2(N263), .B1(n529), .B2(\regOut[10][3] ), .ZN(
        n535) );
  INV_X1 U766 ( .A(n536), .ZN(\regIn[10][2] ) );
  AOI22_X1 U767 ( .A1(n1257), .A2(N263), .B1(n529), .B2(\regOut[10][2] ), .ZN(
        n536) );
  INV_X1 U768 ( .A(n537), .ZN(\regIn[10][1] ) );
  AOI22_X1 U769 ( .A1(n1259), .A2(N263), .B1(n529), .B2(\regOut[10][1] ), .ZN(
        n537) );
  INV_X1 U770 ( .A(n538), .ZN(\regIn[10][15] ) );
  AOI22_X1 U771 ( .A1(n1272), .A2(N263), .B1(n529), .B2(\regOut[10][15] ), 
        .ZN(n538) );
  INV_X1 U772 ( .A(n539), .ZN(\regIn[10][14] ) );
  AOI22_X1 U773 ( .A1(n1270), .A2(N263), .B1(n529), .B2(\regOut[10][14] ), 
        .ZN(n539) );
  INV_X1 U774 ( .A(n540), .ZN(\regIn[10][13] ) );
  AOI22_X1 U775 ( .A1(n1268), .A2(N263), .B1(n529), .B2(\regOut[10][13] ), 
        .ZN(n540) );
  INV_X1 U776 ( .A(n541), .ZN(\regIn[10][12] ) );
  AOI22_X1 U777 ( .A1(n1266), .A2(N263), .B1(n529), .B2(\regOut[10][12] ), 
        .ZN(n541) );
  INV_X1 U778 ( .A(n542), .ZN(\regIn[10][11] ) );
  AOI22_X1 U779 ( .A1(n1264), .A2(N263), .B1(n529), .B2(\regOut[10][11] ), 
        .ZN(n542) );
  INV_X1 U780 ( .A(n543), .ZN(\regIn[10][10] ) );
  AOI22_X1 U781 ( .A1(n1262), .A2(N263), .B1(n529), .B2(\regOut[10][10] ), 
        .ZN(n543) );
  INV_X1 U782 ( .A(n544), .ZN(\regIn[10][0] ) );
  AOI22_X1 U783 ( .A1(n1261), .A2(N263), .B1(n529), .B2(\regOut[10][0] ), .ZN(
        n544) );
  INV_X1 U784 ( .A(N263), .ZN(n529) );
  OAI22_X1 U785 ( .A1(n3), .A2(n545), .B1(N199), .B2(n546), .ZN(\regIn[0][9] )
         );
  INV_X1 U786 ( .A(n1260), .ZN(n3) );
  OAI22_X1 U787 ( .A1(n5), .A2(n545), .B1(N199), .B2(n547), .ZN(\regIn[0][8] )
         );
  INV_X1 U788 ( .A(n1258), .ZN(n5) );
  OAI22_X1 U789 ( .A1(n7), .A2(n545), .B1(N199), .B2(n548), .ZN(\regIn[0][7] )
         );
  INV_X1 U790 ( .A(n1256), .ZN(n7) );
  OAI22_X1 U791 ( .A1(n9), .A2(n545), .B1(N199), .B2(n549), .ZN(\regIn[0][6] )
         );
  INV_X1 U792 ( .A(n1254), .ZN(n9) );
  OAI22_X1 U793 ( .A1(n11), .A2(n545), .B1(N199), .B2(n550), .ZN(\regIn[0][5] ) );
  INV_X1 U794 ( .A(n1252), .ZN(n11) );
  OAI22_X1 U795 ( .A1(n13), .A2(n545), .B1(N199), .B2(n551), .ZN(\regIn[0][4] ) );
  INV_X1 U796 ( .A(n1253), .ZN(n13) );
  OAI22_X1 U797 ( .A1(n15), .A2(n545), .B1(N199), .B2(n552), .ZN(\regIn[0][3] ) );
  INV_X1 U798 ( .A(n1255), .ZN(n15) );
  OAI22_X1 U799 ( .A1(n17), .A2(n545), .B1(N199), .B2(n553), .ZN(\regIn[0][2] ) );
  INV_X1 U800 ( .A(n1257), .ZN(n17) );
  OAI22_X1 U801 ( .A1(n19), .A2(n545), .B1(N199), .B2(n554), .ZN(\regIn[0][1] ) );
  INV_X1 U802 ( .A(n1259), .ZN(n19) );
  OAI22_X1 U803 ( .A1(n21), .A2(n545), .B1(N199), .B2(n555), .ZN(
        \regIn[0][15] ) );
  INV_X1 U804 ( .A(n1272), .ZN(n21) );
  OAI22_X1 U805 ( .A1(n23), .A2(n545), .B1(N199), .B2(n556), .ZN(
        \regIn[0][14] ) );
  INV_X1 U806 ( .A(n1270), .ZN(n23) );
  OAI22_X1 U807 ( .A1(n25), .A2(n545), .B1(N199), .B2(n557), .ZN(
        \regIn[0][13] ) );
  INV_X1 U808 ( .A(n1268), .ZN(n25) );
  OAI22_X1 U809 ( .A1(n27), .A2(n545), .B1(N199), .B2(n558), .ZN(
        \regIn[0][12] ) );
  INV_X1 U810 ( .A(n1266), .ZN(n27) );
  OAI22_X1 U811 ( .A1(n29), .A2(n545), .B1(N199), .B2(n559), .ZN(
        \regIn[0][11] ) );
  INV_X1 U812 ( .A(n1264), .ZN(n29) );
  OAI22_X1 U813 ( .A1(n31), .A2(n545), .B1(N199), .B2(n560), .ZN(
        \regIn[0][10] ) );
  INV_X1 U814 ( .A(n1262), .ZN(n31) );
  OAI22_X1 U815 ( .A1(n33), .A2(n545), .B1(N199), .B2(n561), .ZN(\regIn[0][0] ) );
  INV_X1 U816 ( .A(N199), .ZN(n545) );
  INV_X1 U817 ( .A(n1261), .ZN(n33) );
  NAND2_X1 U818 ( .A1(n562), .A2(n563), .ZN(outB[9]) );
  NOR4_X1 U819 ( .A1(n564), .A2(n565), .A3(n566), .A4(n567), .ZN(n563) );
  OAI221_X1 U820 ( .B1(n410), .B2(n568), .C1(n427), .C2(n569), .A(n570), .ZN(
        n567) );
  AOI22_X1 U821 ( .A1(n571), .A2(\regOut[19][9] ), .B1(n572), .B2(
        \regOut[18][9] ), .ZN(n570) );
  OAI221_X1 U822 ( .B1(n325), .B2(n573), .C1(n342), .C2(n574), .A(n575), .ZN(
        n566) );
  AOI22_X1 U823 ( .A1(n576), .A2(\regOut[23][9] ), .B1(n577), .B2(
        \regOut[22][9] ), .ZN(n575) );
  OAI221_X1 U824 ( .B1(n257), .B2(n578), .C1(n274), .C2(n579), .A(n580), .ZN(
        n565) );
  AOI22_X1 U825 ( .A1(n581), .A2(\regOut[27][9] ), .B1(n582), .B2(
        \regOut[26][9] ), .ZN(n580) );
  OAI221_X1 U826 ( .B1(n138), .B2(n583), .C1(n155), .C2(n584), .A(n585), .ZN(
        n564) );
  AOI22_X1 U827 ( .A1(n586), .A2(\regOut[29][9] ), .B1(n587), .B2(
        \regOut[28][9] ), .ZN(n585) );
  NOR4_X1 U828 ( .A1(n588), .A2(n589), .A3(n590), .A4(n591), .ZN(n562) );
  OAI221_X1 U829 ( .B1(n359), .B2(n592), .C1(n546), .C2(n593), .A(n594), .ZN(
        n591) );
  AOI22_X1 U830 ( .A1(n595), .A2(\regOut[3][9] ), .B1(n596), .B2(
        \regOut[2][9] ), .ZN(n594) );
  OAI221_X1 U831 ( .B1(n87), .B2(n597), .C1(n104), .C2(n598), .A(n599), .ZN(
        n590) );
  AOI22_X1 U832 ( .A1(n600), .A2(\regOut[7][9] ), .B1(n601), .B2(
        \regOut[6][9] ), .ZN(n599) );
  OAI221_X1 U833 ( .B1(n4), .B2(n602), .C1(n36), .C2(n603), .A(n604), .ZN(n589) );
  AOI22_X1 U834 ( .A1(n605), .A2(\regOut[11][9] ), .B1(n606), .B2(
        \regOut[10][9] ), .ZN(n604) );
  OAI221_X1 U835 ( .B1(n478), .B2(n607), .C1(n495), .C2(n608), .A(n609), .ZN(
        n588) );
  AOI22_X1 U836 ( .A1(n610), .A2(\regOut[15][9] ), .B1(n611), .B2(
        \regOut[14][9] ), .ZN(n609) );
  NAND2_X1 U837 ( .A1(n612), .A2(n613), .ZN(outB[8]) );
  NOR4_X1 U838 ( .A1(n614), .A2(n615), .A3(n616), .A4(n617), .ZN(n613) );
  OAI221_X1 U839 ( .B1(n411), .B2(n568), .C1(n428), .C2(n569), .A(n618), .ZN(
        n617) );
  AOI22_X1 U840 ( .A1(n571), .A2(\regOut[19][8] ), .B1(n572), .B2(
        \regOut[18][8] ), .ZN(n618) );
  OAI221_X1 U841 ( .B1(n326), .B2(n573), .C1(n343), .C2(n574), .A(n619), .ZN(
        n616) );
  AOI22_X1 U842 ( .A1(n576), .A2(\regOut[23][8] ), .B1(n577), .B2(
        \regOut[22][8] ), .ZN(n619) );
  OAI221_X1 U843 ( .B1(n258), .B2(n578), .C1(n275), .C2(n579), .A(n620), .ZN(
        n615) );
  AOI22_X1 U844 ( .A1(n581), .A2(\regOut[27][8] ), .B1(n582), .B2(
        \regOut[26][8] ), .ZN(n620) );
  OAI221_X1 U845 ( .B1(n139), .B2(n583), .C1(n156), .C2(n584), .A(n621), .ZN(
        n614) );
  AOI22_X1 U846 ( .A1(n586), .A2(\regOut[29][8] ), .B1(n587), .B2(
        \regOut[28][8] ), .ZN(n621) );
  NOR4_X1 U847 ( .A1(n622), .A2(n623), .A3(n624), .A4(n625), .ZN(n612) );
  OAI221_X1 U848 ( .B1(n360), .B2(n592), .C1(n547), .C2(n593), .A(n626), .ZN(
        n625) );
  AOI22_X1 U849 ( .A1(n595), .A2(\regOut[3][8] ), .B1(n596), .B2(
        \regOut[2][8] ), .ZN(n626) );
  OAI221_X1 U850 ( .B1(n88), .B2(n597), .C1(n105), .C2(n598), .A(n627), .ZN(
        n624) );
  AOI22_X1 U851 ( .A1(n600), .A2(\regOut[7][8] ), .B1(n601), .B2(
        \regOut[6][8] ), .ZN(n627) );
  OAI221_X1 U852 ( .B1(n6), .B2(n602), .C1(n37), .C2(n603), .A(n628), .ZN(n623) );
  AOI22_X1 U853 ( .A1(n605), .A2(\regOut[11][8] ), .B1(n606), .B2(
        \regOut[10][8] ), .ZN(n628) );
  OAI221_X1 U854 ( .B1(n479), .B2(n607), .C1(n496), .C2(n608), .A(n629), .ZN(
        n622) );
  AOI22_X1 U855 ( .A1(n610), .A2(\regOut[15][8] ), .B1(n611), .B2(
        \regOut[14][8] ), .ZN(n629) );
  NAND2_X1 U856 ( .A1(n630), .A2(n631), .ZN(outB[7]) );
  NOR4_X1 U857 ( .A1(n632), .A2(n633), .A3(n634), .A4(n635), .ZN(n631) );
  OAI221_X1 U858 ( .B1(n412), .B2(n568), .C1(n429), .C2(n569), .A(n636), .ZN(
        n635) );
  AOI22_X1 U859 ( .A1(n571), .A2(\regOut[19][7] ), .B1(n572), .B2(
        \regOut[18][7] ), .ZN(n636) );
  OAI221_X1 U860 ( .B1(n327), .B2(n573), .C1(n344), .C2(n574), .A(n637), .ZN(
        n634) );
  AOI22_X1 U861 ( .A1(n576), .A2(\regOut[23][7] ), .B1(n577), .B2(
        \regOut[22][7] ), .ZN(n637) );
  OAI221_X1 U862 ( .B1(n259), .B2(n578), .C1(n276), .C2(n579), .A(n638), .ZN(
        n633) );
  AOI22_X1 U863 ( .A1(n581), .A2(\regOut[27][7] ), .B1(n582), .B2(
        \regOut[26][7] ), .ZN(n638) );
  OAI221_X1 U864 ( .B1(n140), .B2(n583), .C1(n157), .C2(n584), .A(n639), .ZN(
        n632) );
  AOI22_X1 U865 ( .A1(n586), .A2(\regOut[29][7] ), .B1(n587), .B2(
        \regOut[28][7] ), .ZN(n639) );
  NOR4_X1 U866 ( .A1(n640), .A2(n641), .A3(n642), .A4(n643), .ZN(n630) );
  OAI221_X1 U867 ( .B1(n361), .B2(n592), .C1(n548), .C2(n593), .A(n644), .ZN(
        n643) );
  AOI22_X1 U868 ( .A1(n595), .A2(\regOut[3][7] ), .B1(n596), .B2(
        \regOut[2][7] ), .ZN(n644) );
  OAI221_X1 U869 ( .B1(n89), .B2(n597), .C1(n106), .C2(n598), .A(n645), .ZN(
        n642) );
  AOI22_X1 U870 ( .A1(n600), .A2(\regOut[7][7] ), .B1(n601), .B2(
        \regOut[6][7] ), .ZN(n645) );
  OAI221_X1 U871 ( .B1(n8), .B2(n602), .C1(n38), .C2(n603), .A(n646), .ZN(n641) );
  AOI22_X1 U872 ( .A1(n605), .A2(\regOut[11][7] ), .B1(n606), .B2(
        \regOut[10][7] ), .ZN(n646) );
  OAI221_X1 U873 ( .B1(n480), .B2(n607), .C1(n497), .C2(n608), .A(n647), .ZN(
        n640) );
  AOI22_X1 U874 ( .A1(n610), .A2(\regOut[15][7] ), .B1(n611), .B2(
        \regOut[14][7] ), .ZN(n647) );
  NAND2_X1 U875 ( .A1(n648), .A2(n649), .ZN(outB[6]) );
  NOR4_X1 U876 ( .A1(n650), .A2(n651), .A3(n652), .A4(n653), .ZN(n649) );
  OAI221_X1 U877 ( .B1(n413), .B2(n568), .C1(n430), .C2(n569), .A(n654), .ZN(
        n653) );
  AOI22_X1 U878 ( .A1(n571), .A2(\regOut[19][6] ), .B1(n572), .B2(
        \regOut[18][6] ), .ZN(n654) );
  OAI221_X1 U879 ( .B1(n328), .B2(n573), .C1(n345), .C2(n574), .A(n655), .ZN(
        n652) );
  AOI22_X1 U880 ( .A1(n576), .A2(\regOut[23][6] ), .B1(n577), .B2(
        \regOut[22][6] ), .ZN(n655) );
  OAI221_X1 U881 ( .B1(n260), .B2(n578), .C1(n277), .C2(n579), .A(n656), .ZN(
        n651) );
  AOI22_X1 U882 ( .A1(n581), .A2(\regOut[27][6] ), .B1(n582), .B2(
        \regOut[26][6] ), .ZN(n656) );
  OAI221_X1 U883 ( .B1(n141), .B2(n583), .C1(n158), .C2(n584), .A(n657), .ZN(
        n650) );
  AOI22_X1 U884 ( .A1(n586), .A2(\regOut[29][6] ), .B1(n587), .B2(
        \regOut[28][6] ), .ZN(n657) );
  NOR4_X1 U885 ( .A1(n658), .A2(n659), .A3(n660), .A4(n661), .ZN(n648) );
  OAI221_X1 U886 ( .B1(n362), .B2(n592), .C1(n549), .C2(n593), .A(n662), .ZN(
        n661) );
  AOI22_X1 U887 ( .A1(n595), .A2(\regOut[3][6] ), .B1(n596), .B2(
        \regOut[2][6] ), .ZN(n662) );
  OAI221_X1 U888 ( .B1(n90), .B2(n597), .C1(n107), .C2(n598), .A(n663), .ZN(
        n660) );
  AOI22_X1 U889 ( .A1(n600), .A2(\regOut[7][6] ), .B1(n601), .B2(
        \regOut[6][6] ), .ZN(n663) );
  OAI221_X1 U890 ( .B1(n10), .B2(n602), .C1(n39), .C2(n603), .A(n664), .ZN(
        n659) );
  AOI22_X1 U891 ( .A1(n605), .A2(\regOut[11][6] ), .B1(n606), .B2(
        \regOut[10][6] ), .ZN(n664) );
  OAI221_X1 U892 ( .B1(n481), .B2(n607), .C1(n498), .C2(n608), .A(n665), .ZN(
        n658) );
  AOI22_X1 U893 ( .A1(n610), .A2(\regOut[15][6] ), .B1(n611), .B2(
        \regOut[14][6] ), .ZN(n665) );
  NAND2_X1 U894 ( .A1(n666), .A2(n667), .ZN(outB[5]) );
  NOR4_X1 U895 ( .A1(n668), .A2(n669), .A3(n670), .A4(n671), .ZN(n667) );
  OAI221_X1 U896 ( .B1(n414), .B2(n568), .C1(n431), .C2(n569), .A(n672), .ZN(
        n671) );
  AOI22_X1 U897 ( .A1(n571), .A2(\regOut[19][5] ), .B1(n572), .B2(
        \regOut[18][5] ), .ZN(n672) );
  OAI221_X1 U898 ( .B1(n329), .B2(n573), .C1(n346), .C2(n574), .A(n673), .ZN(
        n670) );
  AOI22_X1 U899 ( .A1(n576), .A2(\regOut[23][5] ), .B1(n577), .B2(
        \regOut[22][5] ), .ZN(n673) );
  OAI221_X1 U900 ( .B1(n261), .B2(n578), .C1(n278), .C2(n579), .A(n674), .ZN(
        n669) );
  AOI22_X1 U901 ( .A1(n581), .A2(\regOut[27][5] ), .B1(n582), .B2(
        \regOut[26][5] ), .ZN(n674) );
  OAI221_X1 U902 ( .B1(n142), .B2(n583), .C1(n159), .C2(n584), .A(n675), .ZN(
        n668) );
  AOI22_X1 U903 ( .A1(n586), .A2(\regOut[29][5] ), .B1(n587), .B2(
        \regOut[28][5] ), .ZN(n675) );
  NOR4_X1 U904 ( .A1(n676), .A2(n677), .A3(n678), .A4(n679), .ZN(n666) );
  OAI221_X1 U905 ( .B1(n363), .B2(n592), .C1(n550), .C2(n593), .A(n680), .ZN(
        n679) );
  AOI22_X1 U906 ( .A1(n595), .A2(\regOut[3][5] ), .B1(n596), .B2(
        \regOut[2][5] ), .ZN(n680) );
  OAI221_X1 U907 ( .B1(n91), .B2(n597), .C1(n108), .C2(n598), .A(n681), .ZN(
        n678) );
  AOI22_X1 U908 ( .A1(n600), .A2(\regOut[7][5] ), .B1(n601), .B2(
        \regOut[6][5] ), .ZN(n681) );
  OAI221_X1 U909 ( .B1(n12), .B2(n602), .C1(n40), .C2(n603), .A(n682), .ZN(
        n677) );
  AOI22_X1 U910 ( .A1(n605), .A2(\regOut[11][5] ), .B1(n606), .B2(
        \regOut[10][5] ), .ZN(n682) );
  OAI221_X1 U911 ( .B1(n482), .B2(n607), .C1(n499), .C2(n608), .A(n683), .ZN(
        n676) );
  AOI22_X1 U912 ( .A1(n610), .A2(\regOut[15][5] ), .B1(n611), .B2(
        \regOut[14][5] ), .ZN(n683) );
  NAND2_X1 U913 ( .A1(n684), .A2(n685), .ZN(outB[4]) );
  NOR4_X1 U914 ( .A1(n686), .A2(n687), .A3(n688), .A4(n689), .ZN(n685) );
  OAI221_X1 U915 ( .B1(n415), .B2(n568), .C1(n432), .C2(n569), .A(n690), .ZN(
        n689) );
  AOI22_X1 U916 ( .A1(n571), .A2(\regOut[19][4] ), .B1(n572), .B2(
        \regOut[18][4] ), .ZN(n690) );
  OAI221_X1 U917 ( .B1(n330), .B2(n573), .C1(n347), .C2(n574), .A(n691), .ZN(
        n688) );
  AOI22_X1 U918 ( .A1(n576), .A2(\regOut[23][4] ), .B1(n577), .B2(
        \regOut[22][4] ), .ZN(n691) );
  OAI221_X1 U919 ( .B1(n262), .B2(n578), .C1(n279), .C2(n579), .A(n692), .ZN(
        n687) );
  AOI22_X1 U920 ( .A1(n581), .A2(\regOut[27][4] ), .B1(n582), .B2(
        \regOut[26][4] ), .ZN(n692) );
  OAI221_X1 U921 ( .B1(n143), .B2(n583), .C1(n160), .C2(n584), .A(n693), .ZN(
        n686) );
  AOI22_X1 U922 ( .A1(n586), .A2(\regOut[29][4] ), .B1(n587), .B2(
        \regOut[28][4] ), .ZN(n693) );
  NOR4_X1 U923 ( .A1(n694), .A2(n695), .A3(n696), .A4(n697), .ZN(n684) );
  OAI221_X1 U924 ( .B1(n364), .B2(n592), .C1(n551), .C2(n593), .A(n698), .ZN(
        n697) );
  AOI22_X1 U925 ( .A1(n595), .A2(\regOut[3][4] ), .B1(n596), .B2(
        \regOut[2][4] ), .ZN(n698) );
  OAI221_X1 U926 ( .B1(n92), .B2(n597), .C1(n109), .C2(n598), .A(n699), .ZN(
        n696) );
  AOI22_X1 U927 ( .A1(n600), .A2(\regOut[7][4] ), .B1(n601), .B2(
        \regOut[6][4] ), .ZN(n699) );
  OAI221_X1 U928 ( .B1(n14), .B2(n602), .C1(n41), .C2(n603), .A(n700), .ZN(
        n695) );
  AOI22_X1 U929 ( .A1(n605), .A2(\regOut[11][4] ), .B1(n606), .B2(
        \regOut[10][4] ), .ZN(n700) );
  OAI221_X1 U930 ( .B1(n483), .B2(n607), .C1(n500), .C2(n608), .A(n701), .ZN(
        n694) );
  AOI22_X1 U931 ( .A1(n610), .A2(\regOut[15][4] ), .B1(n611), .B2(
        \regOut[14][4] ), .ZN(n701) );
  NAND2_X1 U932 ( .A1(n702), .A2(n703), .ZN(outB[3]) );
  NOR4_X1 U933 ( .A1(n704), .A2(n705), .A3(n706), .A4(n707), .ZN(n703) );
  OAI221_X1 U934 ( .B1(n416), .B2(n568), .C1(n433), .C2(n569), .A(n708), .ZN(
        n707) );
  AOI22_X1 U935 ( .A1(n571), .A2(\regOut[19][3] ), .B1(n572), .B2(
        \regOut[18][3] ), .ZN(n708) );
  OAI221_X1 U936 ( .B1(n331), .B2(n573), .C1(n348), .C2(n574), .A(n709), .ZN(
        n706) );
  AOI22_X1 U937 ( .A1(n576), .A2(\regOut[23][3] ), .B1(n577), .B2(
        \regOut[22][3] ), .ZN(n709) );
  OAI221_X1 U938 ( .B1(n263), .B2(n578), .C1(n280), .C2(n579), .A(n710), .ZN(
        n705) );
  AOI22_X1 U939 ( .A1(n581), .A2(\regOut[27][3] ), .B1(n582), .B2(
        \regOut[26][3] ), .ZN(n710) );
  OAI221_X1 U940 ( .B1(n144), .B2(n583), .C1(n161), .C2(n584), .A(n711), .ZN(
        n704) );
  AOI22_X1 U941 ( .A1(n586), .A2(\regOut[29][3] ), .B1(n587), .B2(
        \regOut[28][3] ), .ZN(n711) );
  NOR4_X1 U942 ( .A1(n712), .A2(n713), .A3(n714), .A4(n715), .ZN(n702) );
  OAI221_X1 U943 ( .B1(n365), .B2(n592), .C1(n552), .C2(n593), .A(n716), .ZN(
        n715) );
  AOI22_X1 U944 ( .A1(n595), .A2(\regOut[3][3] ), .B1(n596), .B2(
        \regOut[2][3] ), .ZN(n716) );
  OAI221_X1 U945 ( .B1(n93), .B2(n597), .C1(n110), .C2(n598), .A(n717), .ZN(
        n714) );
  AOI22_X1 U946 ( .A1(n600), .A2(\regOut[7][3] ), .B1(n601), .B2(
        \regOut[6][3] ), .ZN(n717) );
  OAI221_X1 U947 ( .B1(n16), .B2(n602), .C1(n42), .C2(n603), .A(n718), .ZN(
        n713) );
  AOI22_X1 U948 ( .A1(n605), .A2(\regOut[11][3] ), .B1(n606), .B2(
        \regOut[10][3] ), .ZN(n718) );
  OAI221_X1 U949 ( .B1(n484), .B2(n607), .C1(n501), .C2(n608), .A(n719), .ZN(
        n712) );
  AOI22_X1 U950 ( .A1(n610), .A2(\regOut[15][3] ), .B1(n611), .B2(
        \regOut[14][3] ), .ZN(n719) );
  NAND2_X1 U951 ( .A1(n720), .A2(n721), .ZN(outB[2]) );
  NOR4_X1 U952 ( .A1(n722), .A2(n723), .A3(n724), .A4(n725), .ZN(n721) );
  OAI221_X1 U953 ( .B1(n417), .B2(n568), .C1(n434), .C2(n569), .A(n726), .ZN(
        n725) );
  AOI22_X1 U954 ( .A1(n571), .A2(\regOut[19][2] ), .B1(n572), .B2(
        \regOut[18][2] ), .ZN(n726) );
  OAI221_X1 U955 ( .B1(n332), .B2(n573), .C1(n349), .C2(n574), .A(n727), .ZN(
        n724) );
  AOI22_X1 U956 ( .A1(n576), .A2(\regOut[23][2] ), .B1(n577), .B2(
        \regOut[22][2] ), .ZN(n727) );
  OAI221_X1 U957 ( .B1(n264), .B2(n578), .C1(n281), .C2(n579), .A(n728), .ZN(
        n723) );
  AOI22_X1 U958 ( .A1(n581), .A2(\regOut[27][2] ), .B1(n582), .B2(
        \regOut[26][2] ), .ZN(n728) );
  OAI221_X1 U959 ( .B1(n145), .B2(n583), .C1(n162), .C2(n584), .A(n729), .ZN(
        n722) );
  AOI22_X1 U960 ( .A1(n586), .A2(\regOut[29][2] ), .B1(n587), .B2(
        \regOut[28][2] ), .ZN(n729) );
  NOR4_X1 U961 ( .A1(n730), .A2(n731), .A3(n732), .A4(n733), .ZN(n720) );
  OAI221_X1 U962 ( .B1(n366), .B2(n592), .C1(n553), .C2(n593), .A(n734), .ZN(
        n733) );
  AOI22_X1 U963 ( .A1(n595), .A2(\regOut[3][2] ), .B1(n596), .B2(
        \regOut[2][2] ), .ZN(n734) );
  OAI221_X1 U964 ( .B1(n94), .B2(n597), .C1(n111), .C2(n598), .A(n735), .ZN(
        n732) );
  AOI22_X1 U965 ( .A1(n600), .A2(\regOut[7][2] ), .B1(n601), .B2(
        \regOut[6][2] ), .ZN(n735) );
  OAI221_X1 U966 ( .B1(n18), .B2(n602), .C1(n43), .C2(n603), .A(n736), .ZN(
        n731) );
  AOI22_X1 U967 ( .A1(n605), .A2(\regOut[11][2] ), .B1(n606), .B2(
        \regOut[10][2] ), .ZN(n736) );
  OAI221_X1 U968 ( .B1(n485), .B2(n607), .C1(n502), .C2(n608), .A(n737), .ZN(
        n730) );
  AOI22_X1 U969 ( .A1(n610), .A2(\regOut[15][2] ), .B1(n611), .B2(
        \regOut[14][2] ), .ZN(n737) );
  NAND2_X1 U970 ( .A1(n738), .A2(n739), .ZN(outB[1]) );
  NOR4_X1 U971 ( .A1(n740), .A2(n741), .A3(n742), .A4(n743), .ZN(n739) );
  OAI221_X1 U972 ( .B1(n418), .B2(n568), .C1(n435), .C2(n569), .A(n744), .ZN(
        n743) );
  AOI22_X1 U973 ( .A1(n571), .A2(\regOut[19][1] ), .B1(n572), .B2(
        \regOut[18][1] ), .ZN(n744) );
  OAI221_X1 U974 ( .B1(n333), .B2(n573), .C1(n350), .C2(n574), .A(n745), .ZN(
        n742) );
  AOI22_X1 U975 ( .A1(n576), .A2(\regOut[23][1] ), .B1(n577), .B2(
        \regOut[22][1] ), .ZN(n745) );
  OAI221_X1 U976 ( .B1(n265), .B2(n578), .C1(n282), .C2(n579), .A(n746), .ZN(
        n741) );
  AOI22_X1 U977 ( .A1(n581), .A2(\regOut[27][1] ), .B1(n582), .B2(
        \regOut[26][1] ), .ZN(n746) );
  OAI221_X1 U978 ( .B1(n146), .B2(n583), .C1(n163), .C2(n584), .A(n747), .ZN(
        n740) );
  AOI22_X1 U979 ( .A1(n586), .A2(\regOut[29][1] ), .B1(n587), .B2(
        \regOut[28][1] ), .ZN(n747) );
  NOR4_X1 U980 ( .A1(n748), .A2(n749), .A3(n750), .A4(n751), .ZN(n738) );
  OAI221_X1 U981 ( .B1(n367), .B2(n592), .C1(n554), .C2(n593), .A(n752), .ZN(
        n751) );
  AOI22_X1 U982 ( .A1(n595), .A2(\regOut[3][1] ), .B1(n596), .B2(
        \regOut[2][1] ), .ZN(n752) );
  OAI221_X1 U983 ( .B1(n95), .B2(n597), .C1(n112), .C2(n598), .A(n753), .ZN(
        n750) );
  AOI22_X1 U984 ( .A1(n600), .A2(\regOut[7][1] ), .B1(n601), .B2(
        \regOut[6][1] ), .ZN(n753) );
  OAI221_X1 U985 ( .B1(n20), .B2(n602), .C1(n44), .C2(n603), .A(n754), .ZN(
        n749) );
  AOI22_X1 U986 ( .A1(n605), .A2(\regOut[11][1] ), .B1(n606), .B2(
        \regOut[10][1] ), .ZN(n754) );
  OAI221_X1 U987 ( .B1(n486), .B2(n607), .C1(n503), .C2(n608), .A(n755), .ZN(
        n748) );
  AOI22_X1 U988 ( .A1(n610), .A2(\regOut[15][1] ), .B1(n611), .B2(
        \regOut[14][1] ), .ZN(n755) );
  NAND2_X1 U989 ( .A1(n756), .A2(n757), .ZN(outB[15]) );
  NOR4_X1 U990 ( .A1(n758), .A2(n759), .A3(n760), .A4(n761), .ZN(n757) );
  OAI221_X1 U991 ( .B1(n419), .B2(n568), .C1(n436), .C2(n569), .A(n762), .ZN(
        n761) );
  AOI22_X1 U992 ( .A1(n571), .A2(\regOut[19][15] ), .B1(n572), .B2(
        \regOut[18][15] ), .ZN(n762) );
  OAI221_X1 U993 ( .B1(n334), .B2(n573), .C1(n351), .C2(n574), .A(n763), .ZN(
        n760) );
  AOI22_X1 U994 ( .A1(n576), .A2(\regOut[23][15] ), .B1(n577), .B2(
        \regOut[22][15] ), .ZN(n763) );
  OAI221_X1 U995 ( .B1(n266), .B2(n578), .C1(n283), .C2(n579), .A(n764), .ZN(
        n759) );
  AOI22_X1 U996 ( .A1(n581), .A2(\regOut[27][15] ), .B1(n582), .B2(
        \regOut[26][15] ), .ZN(n764) );
  OAI221_X1 U997 ( .B1(n147), .B2(n583), .C1(n164), .C2(n584), .A(n765), .ZN(
        n758) );
  AOI22_X1 U998 ( .A1(n586), .A2(\regOut[29][15] ), .B1(n587), .B2(
        \regOut[28][15] ), .ZN(n765) );
  NOR4_X1 U999 ( .A1(n766), .A2(n767), .A3(n768), .A4(n769), .ZN(n756) );
  OAI221_X1 U1000 ( .B1(n368), .B2(n592), .C1(n555), .C2(n593), .A(n770), .ZN(
        n769) );
  AOI22_X1 U1001 ( .A1(n595), .A2(\regOut[3][15] ), .B1(n596), .B2(
        \regOut[2][15] ), .ZN(n770) );
  OAI221_X1 U1002 ( .B1(n96), .B2(n597), .C1(n113), .C2(n598), .A(n771), .ZN(
        n768) );
  AOI22_X1 U1003 ( .A1(n600), .A2(\regOut[7][15] ), .B1(n601), .B2(
        \regOut[6][15] ), .ZN(n771) );
  OAI221_X1 U1004 ( .B1(n22), .B2(n602), .C1(n45), .C2(n603), .A(n772), .ZN(
        n767) );
  AOI22_X1 U1005 ( .A1(n605), .A2(\regOut[11][15] ), .B1(n606), .B2(
        \regOut[10][15] ), .ZN(n772) );
  OAI221_X1 U1006 ( .B1(n487), .B2(n607), .C1(n504), .C2(n608), .A(n773), .ZN(
        n766) );
  AOI22_X1 U1007 ( .A1(n610), .A2(\regOut[15][15] ), .B1(n611), .B2(
        \regOut[14][15] ), .ZN(n773) );
  NAND2_X1 U1008 ( .A1(n774), .A2(n775), .ZN(outB[14]) );
  NOR4_X1 U1009 ( .A1(n776), .A2(n777), .A3(n778), .A4(n779), .ZN(n775) );
  OAI221_X1 U1010 ( .B1(n420), .B2(n568), .C1(n437), .C2(n569), .A(n780), .ZN(
        n779) );
  AOI22_X1 U1011 ( .A1(n571), .A2(\regOut[19][14] ), .B1(n572), .B2(
        \regOut[18][14] ), .ZN(n780) );
  OAI221_X1 U1012 ( .B1(n335), .B2(n573), .C1(n352), .C2(n574), .A(n781), .ZN(
        n778) );
  AOI22_X1 U1013 ( .A1(n576), .A2(\regOut[23][14] ), .B1(n577), .B2(
        \regOut[22][14] ), .ZN(n781) );
  OAI221_X1 U1014 ( .B1(n267), .B2(n578), .C1(n284), .C2(n579), .A(n782), .ZN(
        n777) );
  AOI22_X1 U1015 ( .A1(n581), .A2(\regOut[27][14] ), .B1(n582), .B2(
        \regOut[26][14] ), .ZN(n782) );
  OAI221_X1 U1016 ( .B1(n148), .B2(n583), .C1(n165), .C2(n584), .A(n783), .ZN(
        n776) );
  AOI22_X1 U1017 ( .A1(n586), .A2(\regOut[29][14] ), .B1(n587), .B2(
        \regOut[28][14] ), .ZN(n783) );
  NOR4_X1 U1018 ( .A1(n784), .A2(n785), .A3(n786), .A4(n787), .ZN(n774) );
  OAI221_X1 U1019 ( .B1(n369), .B2(n592), .C1(n556), .C2(n593), .A(n788), .ZN(
        n787) );
  AOI22_X1 U1020 ( .A1(n595), .A2(\regOut[3][14] ), .B1(n596), .B2(
        \regOut[2][14] ), .ZN(n788) );
  OAI221_X1 U1021 ( .B1(n97), .B2(n597), .C1(n114), .C2(n598), .A(n789), .ZN(
        n786) );
  AOI22_X1 U1022 ( .A1(n600), .A2(\regOut[7][14] ), .B1(n601), .B2(
        \regOut[6][14] ), .ZN(n789) );
  OAI221_X1 U1023 ( .B1(n24), .B2(n602), .C1(n46), .C2(n603), .A(n790), .ZN(
        n785) );
  AOI22_X1 U1024 ( .A1(n605), .A2(\regOut[11][14] ), .B1(n606), .B2(
        \regOut[10][14] ), .ZN(n790) );
  OAI221_X1 U1025 ( .B1(n488), .B2(n607), .C1(n505), .C2(n608), .A(n791), .ZN(
        n784) );
  AOI22_X1 U1026 ( .A1(n610), .A2(\regOut[15][14] ), .B1(n611), .B2(
        \regOut[14][14] ), .ZN(n791) );
  NAND2_X1 U1027 ( .A1(n792), .A2(n793), .ZN(outB[13]) );
  NOR4_X1 U1028 ( .A1(n794), .A2(n795), .A3(n796), .A4(n797), .ZN(n793) );
  OAI221_X1 U1029 ( .B1(n421), .B2(n568), .C1(n438), .C2(n569), .A(n798), .ZN(
        n797) );
  AOI22_X1 U1030 ( .A1(n571), .A2(\regOut[19][13] ), .B1(n572), .B2(
        \regOut[18][13] ), .ZN(n798) );
  OAI221_X1 U1031 ( .B1(n336), .B2(n573), .C1(n353), .C2(n574), .A(n799), .ZN(
        n796) );
  AOI22_X1 U1032 ( .A1(n576), .A2(\regOut[23][13] ), .B1(n577), .B2(
        \regOut[22][13] ), .ZN(n799) );
  OAI221_X1 U1033 ( .B1(n268), .B2(n578), .C1(n285), .C2(n579), .A(n800), .ZN(
        n795) );
  AOI22_X1 U1034 ( .A1(n581), .A2(\regOut[27][13] ), .B1(n582), .B2(
        \regOut[26][13] ), .ZN(n800) );
  OAI221_X1 U1035 ( .B1(n149), .B2(n583), .C1(n166), .C2(n584), .A(n801), .ZN(
        n794) );
  AOI22_X1 U1036 ( .A1(n586), .A2(\regOut[29][13] ), .B1(n587), .B2(
        \regOut[28][13] ), .ZN(n801) );
  NOR4_X1 U1037 ( .A1(n802), .A2(n803), .A3(n804), .A4(n805), .ZN(n792) );
  OAI221_X1 U1038 ( .B1(n370), .B2(n592), .C1(n557), .C2(n593), .A(n806), .ZN(
        n805) );
  AOI22_X1 U1039 ( .A1(n595), .A2(\regOut[3][13] ), .B1(n596), .B2(
        \regOut[2][13] ), .ZN(n806) );
  OAI221_X1 U1040 ( .B1(n98), .B2(n597), .C1(n115), .C2(n598), .A(n807), .ZN(
        n804) );
  AOI22_X1 U1041 ( .A1(n600), .A2(\regOut[7][13] ), .B1(n601), .B2(
        \regOut[6][13] ), .ZN(n807) );
  OAI221_X1 U1042 ( .B1(n26), .B2(n602), .C1(n47), .C2(n603), .A(n808), .ZN(
        n803) );
  AOI22_X1 U1043 ( .A1(n605), .A2(\regOut[11][13] ), .B1(n606), .B2(
        \regOut[10][13] ), .ZN(n808) );
  OAI221_X1 U1044 ( .B1(n489), .B2(n607), .C1(n506), .C2(n608), .A(n809), .ZN(
        n802) );
  AOI22_X1 U1045 ( .A1(n610), .A2(\regOut[15][13] ), .B1(n611), .B2(
        \regOut[14][13] ), .ZN(n809) );
  NAND2_X1 U1046 ( .A1(n810), .A2(n811), .ZN(outB[12]) );
  NOR4_X1 U1047 ( .A1(n812), .A2(n813), .A3(n814), .A4(n815), .ZN(n811) );
  OAI221_X1 U1048 ( .B1(n422), .B2(n568), .C1(n439), .C2(n569), .A(n816), .ZN(
        n815) );
  AOI22_X1 U1049 ( .A1(n571), .A2(\regOut[19][12] ), .B1(n572), .B2(
        \regOut[18][12] ), .ZN(n816) );
  OAI221_X1 U1050 ( .B1(n337), .B2(n573), .C1(n354), .C2(n574), .A(n817), .ZN(
        n814) );
  AOI22_X1 U1051 ( .A1(n576), .A2(\regOut[23][12] ), .B1(n577), .B2(
        \regOut[22][12] ), .ZN(n817) );
  OAI221_X1 U1052 ( .B1(n269), .B2(n578), .C1(n286), .C2(n579), .A(n818), .ZN(
        n813) );
  AOI22_X1 U1053 ( .A1(n581), .A2(\regOut[27][12] ), .B1(n582), .B2(
        \regOut[26][12] ), .ZN(n818) );
  OAI221_X1 U1054 ( .B1(n150), .B2(n583), .C1(n167), .C2(n584), .A(n819), .ZN(
        n812) );
  AOI22_X1 U1055 ( .A1(n586), .A2(\regOut[29][12] ), .B1(n587), .B2(
        \regOut[28][12] ), .ZN(n819) );
  NOR4_X1 U1056 ( .A1(n820), .A2(n821), .A3(n822), .A4(n823), .ZN(n810) );
  OAI221_X1 U1057 ( .B1(n371), .B2(n592), .C1(n558), .C2(n593), .A(n824), .ZN(
        n823) );
  AOI22_X1 U1058 ( .A1(n595), .A2(\regOut[3][12] ), .B1(n596), .B2(
        \regOut[2][12] ), .ZN(n824) );
  OAI221_X1 U1059 ( .B1(n99), .B2(n597), .C1(n116), .C2(n598), .A(n825), .ZN(
        n822) );
  AOI22_X1 U1060 ( .A1(n600), .A2(\regOut[7][12] ), .B1(n601), .B2(
        \regOut[6][12] ), .ZN(n825) );
  OAI221_X1 U1061 ( .B1(n28), .B2(n602), .C1(n48), .C2(n603), .A(n826), .ZN(
        n821) );
  AOI22_X1 U1062 ( .A1(n605), .A2(\regOut[11][12] ), .B1(n606), .B2(
        \regOut[10][12] ), .ZN(n826) );
  OAI221_X1 U1063 ( .B1(n490), .B2(n607), .C1(n507), .C2(n608), .A(n827), .ZN(
        n820) );
  AOI22_X1 U1064 ( .A1(n610), .A2(\regOut[15][12] ), .B1(n611), .B2(
        \regOut[14][12] ), .ZN(n827) );
  NAND2_X1 U1065 ( .A1(n828), .A2(n829), .ZN(outB[11]) );
  NOR4_X1 U1066 ( .A1(n830), .A2(n831), .A3(n832), .A4(n833), .ZN(n829) );
  OAI221_X1 U1067 ( .B1(n423), .B2(n568), .C1(n440), .C2(n569), .A(n834), .ZN(
        n833) );
  AOI22_X1 U1068 ( .A1(n571), .A2(\regOut[19][11] ), .B1(n572), .B2(
        \regOut[18][11] ), .ZN(n834) );
  OAI221_X1 U1069 ( .B1(n338), .B2(n573), .C1(n355), .C2(n574), .A(n835), .ZN(
        n832) );
  AOI22_X1 U1070 ( .A1(n576), .A2(\regOut[23][11] ), .B1(n577), .B2(
        \regOut[22][11] ), .ZN(n835) );
  OAI221_X1 U1071 ( .B1(n270), .B2(n578), .C1(n287), .C2(n579), .A(n836), .ZN(
        n831) );
  AOI22_X1 U1072 ( .A1(n581), .A2(\regOut[27][11] ), .B1(n582), .B2(
        \regOut[26][11] ), .ZN(n836) );
  OAI221_X1 U1073 ( .B1(n151), .B2(n583), .C1(n168), .C2(n584), .A(n837), .ZN(
        n830) );
  AOI22_X1 U1074 ( .A1(n586), .A2(\regOut[29][11] ), .B1(n587), .B2(
        \regOut[28][11] ), .ZN(n837) );
  NOR4_X1 U1075 ( .A1(n838), .A2(n839), .A3(n840), .A4(n841), .ZN(n828) );
  OAI221_X1 U1076 ( .B1(n372), .B2(n592), .C1(n559), .C2(n593), .A(n842), .ZN(
        n841) );
  AOI22_X1 U1077 ( .A1(n595), .A2(\regOut[3][11] ), .B1(n596), .B2(
        \regOut[2][11] ), .ZN(n842) );
  OAI221_X1 U1078 ( .B1(n100), .B2(n597), .C1(n117), .C2(n598), .A(n843), .ZN(
        n840) );
  AOI22_X1 U1079 ( .A1(n600), .A2(\regOut[7][11] ), .B1(n601), .B2(
        \regOut[6][11] ), .ZN(n843) );
  OAI221_X1 U1080 ( .B1(n30), .B2(n602), .C1(n49), .C2(n603), .A(n844), .ZN(
        n839) );
  AOI22_X1 U1081 ( .A1(n605), .A2(\regOut[11][11] ), .B1(n606), .B2(
        \regOut[10][11] ), .ZN(n844) );
  OAI221_X1 U1082 ( .B1(n491), .B2(n607), .C1(n508), .C2(n608), .A(n845), .ZN(
        n838) );
  AOI22_X1 U1083 ( .A1(n610), .A2(\regOut[15][11] ), .B1(n611), .B2(
        \regOut[14][11] ), .ZN(n845) );
  NAND2_X1 U1084 ( .A1(n846), .A2(n847), .ZN(outB[10]) );
  NOR4_X1 U1085 ( .A1(n848), .A2(n849), .A3(n850), .A4(n851), .ZN(n847) );
  OAI221_X1 U1086 ( .B1(n424), .B2(n568), .C1(n441), .C2(n569), .A(n852), .ZN(
        n851) );
  AOI22_X1 U1087 ( .A1(n571), .A2(\regOut[19][10] ), .B1(n572), .B2(
        \regOut[18][10] ), .ZN(n852) );
  OAI221_X1 U1088 ( .B1(n339), .B2(n573), .C1(n356), .C2(n574), .A(n853), .ZN(
        n850) );
  AOI22_X1 U1089 ( .A1(n576), .A2(\regOut[23][10] ), .B1(n577), .B2(
        \regOut[22][10] ), .ZN(n853) );
  OAI221_X1 U1090 ( .B1(n271), .B2(n578), .C1(n288), .C2(n579), .A(n854), .ZN(
        n849) );
  AOI22_X1 U1091 ( .A1(n581), .A2(\regOut[27][10] ), .B1(n582), .B2(
        \regOut[26][10] ), .ZN(n854) );
  OAI221_X1 U1092 ( .B1(n152), .B2(n583), .C1(n169), .C2(n584), .A(n855), .ZN(
        n848) );
  AOI22_X1 U1093 ( .A1(n586), .A2(\regOut[29][10] ), .B1(n587), .B2(
        \regOut[28][10] ), .ZN(n855) );
  NOR4_X1 U1094 ( .A1(n856), .A2(n857), .A3(n858), .A4(n859), .ZN(n846) );
  OAI221_X1 U1095 ( .B1(n373), .B2(n592), .C1(n560), .C2(n593), .A(n860), .ZN(
        n859) );
  AOI22_X1 U1096 ( .A1(n595), .A2(\regOut[3][10] ), .B1(n596), .B2(
        \regOut[2][10] ), .ZN(n860) );
  OAI221_X1 U1097 ( .B1(n101), .B2(n597), .C1(n118), .C2(n598), .A(n861), .ZN(
        n858) );
  AOI22_X1 U1098 ( .A1(n600), .A2(\regOut[7][10] ), .B1(n601), .B2(
        \regOut[6][10] ), .ZN(n861) );
  OAI221_X1 U1099 ( .B1(n32), .B2(n602), .C1(n50), .C2(n603), .A(n862), .ZN(
        n857) );
  AOI22_X1 U1100 ( .A1(n605), .A2(\regOut[11][10] ), .B1(n606), .B2(
        \regOut[10][10] ), .ZN(n862) );
  OAI221_X1 U1101 ( .B1(n492), .B2(n607), .C1(n509), .C2(n608), .A(n863), .ZN(
        n856) );
  AOI22_X1 U1102 ( .A1(n610), .A2(\regOut[15][10] ), .B1(n611), .B2(
        \regOut[14][10] ), .ZN(n863) );
  NAND2_X1 U1103 ( .A1(n864), .A2(n865), .ZN(outB[0]) );
  NOR4_X1 U1104 ( .A1(n866), .A2(n867), .A3(n868), .A4(n869), .ZN(n865) );
  OAI221_X1 U1105 ( .B1(n425), .B2(n568), .C1(n442), .C2(n569), .A(n870), .ZN(
        n869) );
  AOI22_X1 U1106 ( .A1(n571), .A2(\regOut[19][0] ), .B1(n572), .B2(
        \regOut[18][0] ), .ZN(n870) );
  AND2_X1 U1107 ( .A1(n871), .A2(n872), .ZN(n572) );
  AND2_X1 U1108 ( .A1(n873), .A2(n872), .ZN(n571) );
  NAND2_X1 U1109 ( .A1(n871), .A2(n874), .ZN(n569) );
  NAND2_X1 U1110 ( .A1(n873), .A2(n874), .ZN(n568) );
  OAI221_X1 U1111 ( .B1(n340), .B2(n573), .C1(n357), .C2(n574), .A(n875), .ZN(
        n868) );
  AOI22_X1 U1112 ( .A1(n576), .A2(\regOut[23][0] ), .B1(n577), .B2(
        \regOut[22][0] ), .ZN(n875) );
  AND2_X1 U1113 ( .A1(n871), .A2(n876), .ZN(n577) );
  AND2_X1 U1114 ( .A1(n873), .A2(n876), .ZN(n576) );
  NAND2_X1 U1115 ( .A1(n871), .A2(n877), .ZN(n574) );
  AND2_X1 U1116 ( .A1(n878), .A2(n879), .ZN(n871) );
  NAND2_X1 U1117 ( .A1(n873), .A2(n877), .ZN(n573) );
  AND2_X1 U1118 ( .A1(n878), .A2(n1251), .ZN(n873) );
  AND2_X1 U1119 ( .A1(n1249), .A2(n880), .ZN(n878) );
  OAI221_X1 U1120 ( .B1(n272), .B2(n578), .C1(n289), .C2(n579), .A(n881), .ZN(
        n867) );
  AOI22_X1 U1121 ( .A1(n581), .A2(\regOut[27][0] ), .B1(n582), .B2(
        \regOut[26][0] ), .ZN(n881) );
  AND2_X1 U1122 ( .A1(n872), .A2(n882), .ZN(n582) );
  AND2_X1 U1123 ( .A1(n872), .A2(n883), .ZN(n581) );
  NAND2_X1 U1124 ( .A1(n874), .A2(n882), .ZN(n579) );
  NAND2_X1 U1125 ( .A1(n874), .A2(n883), .ZN(n578) );
  OAI221_X1 U1126 ( .B1(n153), .B2(n583), .C1(n170), .C2(n584), .A(n884), .ZN(
        n866) );
  AOI22_X1 U1127 ( .A1(n586), .A2(\regOut[29][0] ), .B1(n587), .B2(
        \regOut[28][0] ), .ZN(n884) );
  AND2_X1 U1128 ( .A1(n877), .A2(n882), .ZN(n587) );
  AND2_X1 U1129 ( .A1(n877), .A2(n883), .ZN(n586) );
  NAND2_X1 U1130 ( .A1(n882), .A2(n876), .ZN(n584) );
  AND2_X1 U1131 ( .A1(n885), .A2(n879), .ZN(n882) );
  NAND2_X1 U1132 ( .A1(n876), .A2(n883), .ZN(n583) );
  AND2_X1 U1133 ( .A1(n1251), .A2(n885), .ZN(n883) );
  AND2_X1 U1134 ( .A1(n1249), .A2(n1243), .ZN(n885) );
  NOR4_X1 U1135 ( .A1(n886), .A2(n887), .A3(n888), .A4(n889), .ZN(n864) );
  OAI221_X1 U1136 ( .B1(n374), .B2(n592), .C1(n561), .C2(n593), .A(n890), .ZN(
        n889) );
  AOI22_X1 U1137 ( .A1(n595), .A2(\regOut[3][0] ), .B1(n596), .B2(
        \regOut[2][0] ), .ZN(n890) );
  AND2_X1 U1138 ( .A1(n891), .A2(n872), .ZN(n596) );
  AND2_X1 U1139 ( .A1(n892), .A2(n872), .ZN(n595) );
  NAND2_X1 U1140 ( .A1(n891), .A2(n874), .ZN(n593) );
  NAND2_X1 U1141 ( .A1(n892), .A2(n874), .ZN(n592) );
  OAI221_X1 U1142 ( .B1(n102), .B2(n597), .C1(n119), .C2(n598), .A(n893), .ZN(
        n888) );
  AOI22_X1 U1143 ( .A1(n600), .A2(\regOut[7][0] ), .B1(n601), .B2(
        \regOut[6][0] ), .ZN(n893) );
  AND2_X1 U1144 ( .A1(n891), .A2(n876), .ZN(n601) );
  AND2_X1 U1145 ( .A1(n892), .A2(n876), .ZN(n600) );
  NAND2_X1 U1146 ( .A1(n891), .A2(n877), .ZN(n598) );
  AND2_X1 U1147 ( .A1(n894), .A2(n879), .ZN(n891) );
  NAND2_X1 U1148 ( .A1(n892), .A2(n877), .ZN(n597) );
  AND2_X1 U1149 ( .A1(n894), .A2(n1251), .ZN(n892) );
  NOR2_X1 U1150 ( .A1(n1243), .A2(n1249), .ZN(n894) );
  OAI221_X1 U1151 ( .B1(n34), .B2(n602), .C1(n51), .C2(n603), .A(n895), .ZN(
        n887) );
  AOI22_X1 U1152 ( .A1(n605), .A2(\regOut[11][0] ), .B1(n606), .B2(
        \regOut[10][0] ), .ZN(n895) );
  AND2_X1 U1153 ( .A1(n896), .A2(n872), .ZN(n606) );
  AND2_X1 U1154 ( .A1(n897), .A2(n872), .ZN(n605) );
  NOR2_X1 U1155 ( .A1(n898), .A2(n1245), .ZN(n872) );
  NAND2_X1 U1156 ( .A1(n896), .A2(n874), .ZN(n603) );
  NAND2_X1 U1157 ( .A1(n897), .A2(n874), .ZN(n602) );
  NOR2_X1 U1158 ( .A1(n1247), .A2(n1245), .ZN(n874) );
  OAI221_X1 U1159 ( .B1(n493), .B2(n607), .C1(n510), .C2(n608), .A(n899), .ZN(
        n886) );
  AOI22_X1 U1160 ( .A1(n610), .A2(\regOut[15][0] ), .B1(n611), .B2(
        \regOut[14][0] ), .ZN(n899) );
  AND2_X1 U1161 ( .A1(n896), .A2(n876), .ZN(n611) );
  AND2_X1 U1162 ( .A1(n897), .A2(n876), .ZN(n610) );
  NOR2_X1 U1163 ( .A1(n900), .A2(n898), .ZN(n876) );
  INV_X1 U1164 ( .A(n1247), .ZN(n898) );
  NAND2_X1 U1165 ( .A1(n896), .A2(n877), .ZN(n608) );
  AND2_X1 U1166 ( .A1(n901), .A2(n879), .ZN(n896) );
  INV_X1 U1167 ( .A(n1251), .ZN(n879) );
  NAND2_X1 U1168 ( .A1(n897), .A2(n877), .ZN(n607) );
  NOR2_X1 U1169 ( .A1(n900), .A2(n1247), .ZN(n877) );
  INV_X1 U1170 ( .A(n1245), .ZN(n900) );
  AND2_X1 U1171 ( .A1(n901), .A2(n1251), .ZN(n897) );
  NOR2_X1 U1172 ( .A1(n880), .A2(n1249), .ZN(n901) );
  INV_X1 U1173 ( .A(n1243), .ZN(n880) );
  NAND2_X1 U1174 ( .A1(n902), .A2(n903), .ZN(outA[9]) );
  NOR4_X1 U1175 ( .A1(n904), .A2(n905), .A3(n906), .A4(n907), .ZN(n903) );
  OAI221_X1 U1176 ( .B1(n410), .B2(n908), .C1(n427), .C2(n909), .A(n910), .ZN(
        n907) );
  AOI22_X1 U1177 ( .A1(n911), .A2(\regOut[19][9] ), .B1(n912), .B2(
        \regOut[18][9] ), .ZN(n910) );
  INV_X1 U1178 ( .A(\regOut[16][9] ), .ZN(n427) );
  INV_X1 U1179 ( .A(\regOut[17][9] ), .ZN(n410) );
  OAI221_X1 U1180 ( .B1(n325), .B2(n913), .C1(n342), .C2(n914), .A(n915), .ZN(
        n906) );
  AOI22_X1 U1181 ( .A1(n916), .A2(\regOut[23][9] ), .B1(n917), .B2(
        \regOut[22][9] ), .ZN(n915) );
  INV_X1 U1182 ( .A(\regOut[20][9] ), .ZN(n342) );
  INV_X1 U1183 ( .A(\regOut[21][9] ), .ZN(n325) );
  OAI221_X1 U1184 ( .B1(n257), .B2(n918), .C1(n274), .C2(n919), .A(n920), .ZN(
        n905) );
  AOI22_X1 U1185 ( .A1(n921), .A2(\regOut[27][9] ), .B1(n922), .B2(
        \regOut[26][9] ), .ZN(n920) );
  INV_X1 U1186 ( .A(\regOut[24][9] ), .ZN(n274) );
  INV_X1 U1187 ( .A(\regOut[25][9] ), .ZN(n257) );
  OAI221_X1 U1188 ( .B1(n138), .B2(n923), .C1(n155), .C2(n924), .A(n925), .ZN(
        n904) );
  AOI22_X1 U1189 ( .A1(n926), .A2(\regOut[29][9] ), .B1(n927), .B2(
        \regOut[28][9] ), .ZN(n925) );
  INV_X1 U1190 ( .A(\regOut[30][9] ), .ZN(n155) );
  INV_X1 U1191 ( .A(\regOut[31][9] ), .ZN(n138) );
  NOR4_X1 U1192 ( .A1(n928), .A2(n929), .A3(n930), .A4(n931), .ZN(n902) );
  OAI221_X1 U1193 ( .B1(n359), .B2(n932), .C1(n546), .C2(n933), .A(n934), .ZN(
        n931) );
  AOI22_X1 U1194 ( .A1(n935), .A2(\regOut[3][9] ), .B1(n936), .B2(
        \regOut[2][9] ), .ZN(n934) );
  INV_X1 U1195 ( .A(\regOut[0][9] ), .ZN(n546) );
  INV_X1 U1196 ( .A(\regOut[1][9] ), .ZN(n359) );
  OAI221_X1 U1197 ( .B1(n87), .B2(n937), .C1(n104), .C2(n938), .A(n939), .ZN(
        n930) );
  AOI22_X1 U1198 ( .A1(n940), .A2(\regOut[7][9] ), .B1(n941), .B2(
        \regOut[6][9] ), .ZN(n939) );
  INV_X1 U1199 ( .A(\regOut[4][9] ), .ZN(n104) );
  INV_X1 U1200 ( .A(\regOut[5][9] ), .ZN(n87) );
  OAI221_X1 U1201 ( .B1(n4), .B2(n942), .C1(n36), .C2(n943), .A(n944), .ZN(
        n929) );
  AOI22_X1 U1202 ( .A1(n945), .A2(\regOut[11][9] ), .B1(n946), .B2(
        \regOut[10][9] ), .ZN(n944) );
  INV_X1 U1203 ( .A(\regOut[8][9] ), .ZN(n36) );
  INV_X1 U1204 ( .A(\regOut[9][9] ), .ZN(n4) );
  OAI221_X1 U1205 ( .B1(n478), .B2(n947), .C1(n495), .C2(n948), .A(n949), .ZN(
        n928) );
  AOI22_X1 U1206 ( .A1(n950), .A2(\regOut[15][9] ), .B1(n951), .B2(
        \regOut[14][9] ), .ZN(n949) );
  INV_X1 U1207 ( .A(\regOut[12][9] ), .ZN(n495) );
  INV_X1 U1208 ( .A(\regOut[13][9] ), .ZN(n478) );
  NAND2_X1 U1209 ( .A1(n952), .A2(n953), .ZN(outA[8]) );
  NOR4_X1 U1210 ( .A1(n954), .A2(n955), .A3(n956), .A4(n957), .ZN(n953) );
  OAI221_X1 U1211 ( .B1(n411), .B2(n908), .C1(n428), .C2(n909), .A(n958), .ZN(
        n957) );
  AOI22_X1 U1212 ( .A1(n911), .A2(\regOut[19][8] ), .B1(n912), .B2(
        \regOut[18][8] ), .ZN(n958) );
  INV_X1 U1213 ( .A(\regOut[16][8] ), .ZN(n428) );
  INV_X1 U1214 ( .A(\regOut[17][8] ), .ZN(n411) );
  OAI221_X1 U1215 ( .B1(n326), .B2(n913), .C1(n343), .C2(n914), .A(n959), .ZN(
        n956) );
  AOI22_X1 U1216 ( .A1(n916), .A2(\regOut[23][8] ), .B1(n917), .B2(
        \regOut[22][8] ), .ZN(n959) );
  INV_X1 U1217 ( .A(\regOut[20][8] ), .ZN(n343) );
  INV_X1 U1218 ( .A(\regOut[21][8] ), .ZN(n326) );
  OAI221_X1 U1219 ( .B1(n258), .B2(n918), .C1(n275), .C2(n919), .A(n960), .ZN(
        n955) );
  AOI22_X1 U1220 ( .A1(n921), .A2(\regOut[27][8] ), .B1(n922), .B2(
        \regOut[26][8] ), .ZN(n960) );
  INV_X1 U1221 ( .A(\regOut[24][8] ), .ZN(n275) );
  INV_X1 U1222 ( .A(\regOut[25][8] ), .ZN(n258) );
  OAI221_X1 U1223 ( .B1(n139), .B2(n923), .C1(n156), .C2(n924), .A(n961), .ZN(
        n954) );
  AOI22_X1 U1224 ( .A1(n926), .A2(\regOut[29][8] ), .B1(n927), .B2(
        \regOut[28][8] ), .ZN(n961) );
  INV_X1 U1225 ( .A(\regOut[30][8] ), .ZN(n156) );
  INV_X1 U1226 ( .A(\regOut[31][8] ), .ZN(n139) );
  NOR4_X1 U1227 ( .A1(n962), .A2(n963), .A3(n964), .A4(n965), .ZN(n952) );
  OAI221_X1 U1228 ( .B1(n360), .B2(n932), .C1(n547), .C2(n933), .A(n966), .ZN(
        n965) );
  AOI22_X1 U1229 ( .A1(n935), .A2(\regOut[3][8] ), .B1(n936), .B2(
        \regOut[2][8] ), .ZN(n966) );
  INV_X1 U1230 ( .A(\regOut[0][8] ), .ZN(n547) );
  INV_X1 U1231 ( .A(\regOut[1][8] ), .ZN(n360) );
  OAI221_X1 U1232 ( .B1(n88), .B2(n937), .C1(n105), .C2(n938), .A(n967), .ZN(
        n964) );
  AOI22_X1 U1233 ( .A1(n940), .A2(\regOut[7][8] ), .B1(n941), .B2(
        \regOut[6][8] ), .ZN(n967) );
  INV_X1 U1234 ( .A(\regOut[4][8] ), .ZN(n105) );
  INV_X1 U1235 ( .A(\regOut[5][8] ), .ZN(n88) );
  OAI221_X1 U1236 ( .B1(n6), .B2(n942), .C1(n37), .C2(n943), .A(n968), .ZN(
        n963) );
  AOI22_X1 U1237 ( .A1(n945), .A2(\regOut[11][8] ), .B1(n946), .B2(
        \regOut[10][8] ), .ZN(n968) );
  INV_X1 U1238 ( .A(\regOut[8][8] ), .ZN(n37) );
  INV_X1 U1239 ( .A(\regOut[9][8] ), .ZN(n6) );
  OAI221_X1 U1240 ( .B1(n479), .B2(n947), .C1(n496), .C2(n948), .A(n969), .ZN(
        n962) );
  AOI22_X1 U1241 ( .A1(n950), .A2(\regOut[15][8] ), .B1(n951), .B2(
        \regOut[14][8] ), .ZN(n969) );
  INV_X1 U1242 ( .A(\regOut[12][8] ), .ZN(n496) );
  INV_X1 U1243 ( .A(\regOut[13][8] ), .ZN(n479) );
  NAND2_X1 U1244 ( .A1(n970), .A2(n971), .ZN(outA[7]) );
  NOR4_X1 U1245 ( .A1(n972), .A2(n973), .A3(n974), .A4(n975), .ZN(n971) );
  OAI221_X1 U1246 ( .B1(n412), .B2(n908), .C1(n429), .C2(n909), .A(n976), .ZN(
        n975) );
  AOI22_X1 U1247 ( .A1(n911), .A2(\regOut[19][7] ), .B1(n912), .B2(
        \regOut[18][7] ), .ZN(n976) );
  INV_X1 U1248 ( .A(\regOut[16][7] ), .ZN(n429) );
  INV_X1 U1249 ( .A(\regOut[17][7] ), .ZN(n412) );
  OAI221_X1 U1250 ( .B1(n327), .B2(n913), .C1(n344), .C2(n914), .A(n977), .ZN(
        n974) );
  AOI22_X1 U1251 ( .A1(n916), .A2(\regOut[23][7] ), .B1(n917), .B2(
        \regOut[22][7] ), .ZN(n977) );
  INV_X1 U1252 ( .A(\regOut[20][7] ), .ZN(n344) );
  INV_X1 U1253 ( .A(\regOut[21][7] ), .ZN(n327) );
  OAI221_X1 U1254 ( .B1(n259), .B2(n918), .C1(n276), .C2(n919), .A(n978), .ZN(
        n973) );
  AOI22_X1 U1255 ( .A1(n921), .A2(\regOut[27][7] ), .B1(n922), .B2(
        \regOut[26][7] ), .ZN(n978) );
  INV_X1 U1256 ( .A(\regOut[24][7] ), .ZN(n276) );
  INV_X1 U1257 ( .A(\regOut[25][7] ), .ZN(n259) );
  OAI221_X1 U1258 ( .B1(n140), .B2(n923), .C1(n157), .C2(n924), .A(n979), .ZN(
        n972) );
  AOI22_X1 U1259 ( .A1(n926), .A2(\regOut[29][7] ), .B1(n927), .B2(
        \regOut[28][7] ), .ZN(n979) );
  INV_X1 U1260 ( .A(\regOut[30][7] ), .ZN(n157) );
  INV_X1 U1261 ( .A(\regOut[31][7] ), .ZN(n140) );
  NOR4_X1 U1262 ( .A1(n980), .A2(n981), .A3(n982), .A4(n983), .ZN(n970) );
  OAI221_X1 U1263 ( .B1(n361), .B2(n932), .C1(n548), .C2(n933), .A(n984), .ZN(
        n983) );
  AOI22_X1 U1264 ( .A1(n935), .A2(\regOut[3][7] ), .B1(n936), .B2(
        \regOut[2][7] ), .ZN(n984) );
  INV_X1 U1265 ( .A(\regOut[0][7] ), .ZN(n548) );
  INV_X1 U1266 ( .A(\regOut[1][7] ), .ZN(n361) );
  OAI221_X1 U1267 ( .B1(n89), .B2(n937), .C1(n106), .C2(n938), .A(n985), .ZN(
        n982) );
  AOI22_X1 U1268 ( .A1(n940), .A2(\regOut[7][7] ), .B1(n941), .B2(
        \regOut[6][7] ), .ZN(n985) );
  INV_X1 U1269 ( .A(\regOut[4][7] ), .ZN(n106) );
  INV_X1 U1270 ( .A(\regOut[5][7] ), .ZN(n89) );
  OAI221_X1 U1271 ( .B1(n8), .B2(n942), .C1(n38), .C2(n943), .A(n986), .ZN(
        n981) );
  AOI22_X1 U1272 ( .A1(n945), .A2(\regOut[11][7] ), .B1(n946), .B2(
        \regOut[10][7] ), .ZN(n986) );
  INV_X1 U1273 ( .A(\regOut[8][7] ), .ZN(n38) );
  INV_X1 U1274 ( .A(\regOut[9][7] ), .ZN(n8) );
  OAI221_X1 U1275 ( .B1(n480), .B2(n947), .C1(n497), .C2(n948), .A(n987), .ZN(
        n980) );
  AOI22_X1 U1276 ( .A1(n950), .A2(\regOut[15][7] ), .B1(n951), .B2(
        \regOut[14][7] ), .ZN(n987) );
  INV_X1 U1277 ( .A(\regOut[12][7] ), .ZN(n497) );
  INV_X1 U1278 ( .A(\regOut[13][7] ), .ZN(n480) );
  NAND2_X1 U1279 ( .A1(n988), .A2(n989), .ZN(outA[6]) );
  NOR4_X1 U1280 ( .A1(n990), .A2(n991), .A3(n992), .A4(n993), .ZN(n989) );
  OAI221_X1 U1281 ( .B1(n413), .B2(n908), .C1(n430), .C2(n909), .A(n994), .ZN(
        n993) );
  AOI22_X1 U1282 ( .A1(n911), .A2(\regOut[19][6] ), .B1(n912), .B2(
        \regOut[18][6] ), .ZN(n994) );
  INV_X1 U1283 ( .A(\regOut[16][6] ), .ZN(n430) );
  INV_X1 U1284 ( .A(\regOut[17][6] ), .ZN(n413) );
  OAI221_X1 U1285 ( .B1(n328), .B2(n913), .C1(n345), .C2(n914), .A(n995), .ZN(
        n992) );
  AOI22_X1 U1286 ( .A1(n916), .A2(\regOut[23][6] ), .B1(n917), .B2(
        \regOut[22][6] ), .ZN(n995) );
  INV_X1 U1287 ( .A(\regOut[20][6] ), .ZN(n345) );
  INV_X1 U1288 ( .A(\regOut[21][6] ), .ZN(n328) );
  OAI221_X1 U1289 ( .B1(n260), .B2(n918), .C1(n277), .C2(n919), .A(n996), .ZN(
        n991) );
  AOI22_X1 U1290 ( .A1(n921), .A2(\regOut[27][6] ), .B1(n922), .B2(
        \regOut[26][6] ), .ZN(n996) );
  INV_X1 U1291 ( .A(\regOut[24][6] ), .ZN(n277) );
  INV_X1 U1292 ( .A(\regOut[25][6] ), .ZN(n260) );
  OAI221_X1 U1293 ( .B1(n141), .B2(n923), .C1(n158), .C2(n924), .A(n997), .ZN(
        n990) );
  AOI22_X1 U1294 ( .A1(n926), .A2(\regOut[29][6] ), .B1(n927), .B2(
        \regOut[28][6] ), .ZN(n997) );
  INV_X1 U1295 ( .A(\regOut[30][6] ), .ZN(n158) );
  INV_X1 U1296 ( .A(\regOut[31][6] ), .ZN(n141) );
  NOR4_X1 U1297 ( .A1(n998), .A2(n999), .A3(n1000), .A4(n1001), .ZN(n988) );
  OAI221_X1 U1298 ( .B1(n362), .B2(n932), .C1(n549), .C2(n933), .A(n1002), 
        .ZN(n1001) );
  AOI22_X1 U1299 ( .A1(n935), .A2(\regOut[3][6] ), .B1(n936), .B2(
        \regOut[2][6] ), .ZN(n1002) );
  INV_X1 U1300 ( .A(\regOut[0][6] ), .ZN(n549) );
  INV_X1 U1301 ( .A(\regOut[1][6] ), .ZN(n362) );
  OAI221_X1 U1302 ( .B1(n90), .B2(n937), .C1(n107), .C2(n938), .A(n1003), .ZN(
        n1000) );
  AOI22_X1 U1303 ( .A1(n940), .A2(\regOut[7][6] ), .B1(n941), .B2(
        \regOut[6][6] ), .ZN(n1003) );
  INV_X1 U1304 ( .A(\regOut[4][6] ), .ZN(n107) );
  INV_X1 U1305 ( .A(\regOut[5][6] ), .ZN(n90) );
  OAI221_X1 U1306 ( .B1(n10), .B2(n942), .C1(n39), .C2(n943), .A(n1004), .ZN(
        n999) );
  AOI22_X1 U1307 ( .A1(n945), .A2(\regOut[11][6] ), .B1(n946), .B2(
        \regOut[10][6] ), .ZN(n1004) );
  INV_X1 U1308 ( .A(\regOut[8][6] ), .ZN(n39) );
  INV_X1 U1309 ( .A(\regOut[9][6] ), .ZN(n10) );
  OAI221_X1 U1310 ( .B1(n481), .B2(n947), .C1(n498), .C2(n948), .A(n1005), 
        .ZN(n998) );
  AOI22_X1 U1311 ( .A1(n950), .A2(\regOut[15][6] ), .B1(n951), .B2(
        \regOut[14][6] ), .ZN(n1005) );
  INV_X1 U1312 ( .A(\regOut[12][6] ), .ZN(n498) );
  INV_X1 U1313 ( .A(\regOut[13][6] ), .ZN(n481) );
  NAND2_X1 U1314 ( .A1(n1006), .A2(n1007), .ZN(outA[5]) );
  NOR4_X1 U1315 ( .A1(n1008), .A2(n1009), .A3(n1010), .A4(n1011), .ZN(n1007)
         );
  OAI221_X1 U1316 ( .B1(n414), .B2(n908), .C1(n431), .C2(n909), .A(n1012), 
        .ZN(n1011) );
  AOI22_X1 U1317 ( .A1(n911), .A2(\regOut[19][5] ), .B1(n912), .B2(
        \regOut[18][5] ), .ZN(n1012) );
  INV_X1 U1318 ( .A(\regOut[16][5] ), .ZN(n431) );
  INV_X1 U1319 ( .A(\regOut[17][5] ), .ZN(n414) );
  OAI221_X1 U1320 ( .B1(n329), .B2(n913), .C1(n346), .C2(n914), .A(n1013), 
        .ZN(n1010) );
  AOI22_X1 U1321 ( .A1(n916), .A2(\regOut[23][5] ), .B1(n917), .B2(
        \regOut[22][5] ), .ZN(n1013) );
  INV_X1 U1322 ( .A(\regOut[20][5] ), .ZN(n346) );
  INV_X1 U1323 ( .A(\regOut[21][5] ), .ZN(n329) );
  OAI221_X1 U1324 ( .B1(n261), .B2(n918), .C1(n278), .C2(n919), .A(n1014), 
        .ZN(n1009) );
  AOI22_X1 U1325 ( .A1(n921), .A2(\regOut[27][5] ), .B1(n922), .B2(
        \regOut[26][5] ), .ZN(n1014) );
  INV_X1 U1326 ( .A(\regOut[24][5] ), .ZN(n278) );
  INV_X1 U1327 ( .A(\regOut[25][5] ), .ZN(n261) );
  OAI221_X1 U1328 ( .B1(n142), .B2(n923), .C1(n159), .C2(n924), .A(n1015), 
        .ZN(n1008) );
  AOI22_X1 U1329 ( .A1(n926), .A2(\regOut[29][5] ), .B1(n927), .B2(
        \regOut[28][5] ), .ZN(n1015) );
  INV_X1 U1330 ( .A(\regOut[30][5] ), .ZN(n159) );
  INV_X1 U1331 ( .A(\regOut[31][5] ), .ZN(n142) );
  NOR4_X1 U1332 ( .A1(n1016), .A2(n1017), .A3(n1018), .A4(n1019), .ZN(n1006)
         );
  OAI221_X1 U1333 ( .B1(n363), .B2(n932), .C1(n550), .C2(n933), .A(n1020), 
        .ZN(n1019) );
  AOI22_X1 U1334 ( .A1(n935), .A2(\regOut[3][5] ), .B1(n936), .B2(
        \regOut[2][5] ), .ZN(n1020) );
  INV_X1 U1335 ( .A(\regOut[0][5] ), .ZN(n550) );
  INV_X1 U1336 ( .A(\regOut[1][5] ), .ZN(n363) );
  OAI221_X1 U1337 ( .B1(n91), .B2(n937), .C1(n108), .C2(n938), .A(n1021), .ZN(
        n1018) );
  AOI22_X1 U1338 ( .A1(n940), .A2(\regOut[7][5] ), .B1(n941), .B2(
        \regOut[6][5] ), .ZN(n1021) );
  INV_X1 U1339 ( .A(\regOut[4][5] ), .ZN(n108) );
  INV_X1 U1340 ( .A(\regOut[5][5] ), .ZN(n91) );
  OAI221_X1 U1341 ( .B1(n12), .B2(n942), .C1(n40), .C2(n943), .A(n1022), .ZN(
        n1017) );
  AOI22_X1 U1342 ( .A1(n945), .A2(\regOut[11][5] ), .B1(n946), .B2(
        \regOut[10][5] ), .ZN(n1022) );
  INV_X1 U1343 ( .A(\regOut[8][5] ), .ZN(n40) );
  INV_X1 U1344 ( .A(\regOut[9][5] ), .ZN(n12) );
  OAI221_X1 U1345 ( .B1(n482), .B2(n947), .C1(n499), .C2(n948), .A(n1023), 
        .ZN(n1016) );
  AOI22_X1 U1346 ( .A1(n950), .A2(\regOut[15][5] ), .B1(n951), .B2(
        \regOut[14][5] ), .ZN(n1023) );
  INV_X1 U1347 ( .A(\regOut[12][5] ), .ZN(n499) );
  INV_X1 U1348 ( .A(\regOut[13][5] ), .ZN(n482) );
  NAND2_X1 U1349 ( .A1(n1024), .A2(n1025), .ZN(outA[4]) );
  NOR4_X1 U1350 ( .A1(n1026), .A2(n1027), .A3(n1028), .A4(n1029), .ZN(n1025)
         );
  OAI221_X1 U1351 ( .B1(n415), .B2(n908), .C1(n432), .C2(n909), .A(n1030), 
        .ZN(n1029) );
  AOI22_X1 U1352 ( .A1(n911), .A2(\regOut[19][4] ), .B1(n912), .B2(
        \regOut[18][4] ), .ZN(n1030) );
  INV_X1 U1353 ( .A(\regOut[16][4] ), .ZN(n432) );
  INV_X1 U1354 ( .A(\regOut[17][4] ), .ZN(n415) );
  OAI221_X1 U1355 ( .B1(n330), .B2(n913), .C1(n347), .C2(n914), .A(n1031), 
        .ZN(n1028) );
  AOI22_X1 U1356 ( .A1(n916), .A2(\regOut[23][4] ), .B1(n917), .B2(
        \regOut[22][4] ), .ZN(n1031) );
  INV_X1 U1357 ( .A(\regOut[20][4] ), .ZN(n347) );
  INV_X1 U1358 ( .A(\regOut[21][4] ), .ZN(n330) );
  OAI221_X1 U1359 ( .B1(n262), .B2(n918), .C1(n279), .C2(n919), .A(n1032), 
        .ZN(n1027) );
  AOI22_X1 U1360 ( .A1(n921), .A2(\regOut[27][4] ), .B1(n922), .B2(
        \regOut[26][4] ), .ZN(n1032) );
  INV_X1 U1361 ( .A(\regOut[24][4] ), .ZN(n279) );
  INV_X1 U1362 ( .A(\regOut[25][4] ), .ZN(n262) );
  OAI221_X1 U1363 ( .B1(n143), .B2(n923), .C1(n160), .C2(n924), .A(n1033), 
        .ZN(n1026) );
  AOI22_X1 U1364 ( .A1(n926), .A2(\regOut[29][4] ), .B1(n927), .B2(
        \regOut[28][4] ), .ZN(n1033) );
  INV_X1 U1365 ( .A(\regOut[30][4] ), .ZN(n160) );
  INV_X1 U1366 ( .A(\regOut[31][4] ), .ZN(n143) );
  NOR4_X1 U1367 ( .A1(n1034), .A2(n1035), .A3(n1036), .A4(n1037), .ZN(n1024)
         );
  OAI221_X1 U1368 ( .B1(n364), .B2(n932), .C1(n551), .C2(n933), .A(n1038), 
        .ZN(n1037) );
  AOI22_X1 U1369 ( .A1(n935), .A2(\regOut[3][4] ), .B1(n936), .B2(
        \regOut[2][4] ), .ZN(n1038) );
  INV_X1 U1370 ( .A(\regOut[0][4] ), .ZN(n551) );
  INV_X1 U1371 ( .A(\regOut[1][4] ), .ZN(n364) );
  OAI221_X1 U1372 ( .B1(n92), .B2(n937), .C1(n109), .C2(n938), .A(n1039), .ZN(
        n1036) );
  AOI22_X1 U1373 ( .A1(n940), .A2(\regOut[7][4] ), .B1(n941), .B2(
        \regOut[6][4] ), .ZN(n1039) );
  INV_X1 U1374 ( .A(\regOut[4][4] ), .ZN(n109) );
  INV_X1 U1375 ( .A(\regOut[5][4] ), .ZN(n92) );
  OAI221_X1 U1376 ( .B1(n14), .B2(n942), .C1(n41), .C2(n943), .A(n1040), .ZN(
        n1035) );
  AOI22_X1 U1377 ( .A1(n945), .A2(\regOut[11][4] ), .B1(n946), .B2(
        \regOut[10][4] ), .ZN(n1040) );
  INV_X1 U1378 ( .A(\regOut[8][4] ), .ZN(n41) );
  INV_X1 U1379 ( .A(\regOut[9][4] ), .ZN(n14) );
  OAI221_X1 U1380 ( .B1(n483), .B2(n947), .C1(n500), .C2(n948), .A(n1041), 
        .ZN(n1034) );
  AOI22_X1 U1381 ( .A1(n950), .A2(\regOut[15][4] ), .B1(n951), .B2(
        \regOut[14][4] ), .ZN(n1041) );
  INV_X1 U1382 ( .A(\regOut[12][4] ), .ZN(n500) );
  INV_X1 U1383 ( .A(\regOut[13][4] ), .ZN(n483) );
  NAND2_X1 U1384 ( .A1(n1042), .A2(n1043), .ZN(outA[3]) );
  NOR4_X1 U1385 ( .A1(n1044), .A2(n1045), .A3(n1046), .A4(n1047), .ZN(n1043)
         );
  OAI221_X1 U1386 ( .B1(n416), .B2(n908), .C1(n433), .C2(n909), .A(n1048), 
        .ZN(n1047) );
  AOI22_X1 U1387 ( .A1(n911), .A2(\regOut[19][3] ), .B1(n912), .B2(
        \regOut[18][3] ), .ZN(n1048) );
  INV_X1 U1388 ( .A(\regOut[16][3] ), .ZN(n433) );
  INV_X1 U1389 ( .A(\regOut[17][3] ), .ZN(n416) );
  OAI221_X1 U1390 ( .B1(n331), .B2(n913), .C1(n348), .C2(n914), .A(n1049), 
        .ZN(n1046) );
  AOI22_X1 U1391 ( .A1(n916), .A2(\regOut[23][3] ), .B1(n917), .B2(
        \regOut[22][3] ), .ZN(n1049) );
  INV_X1 U1392 ( .A(\regOut[20][3] ), .ZN(n348) );
  INV_X1 U1393 ( .A(\regOut[21][3] ), .ZN(n331) );
  OAI221_X1 U1394 ( .B1(n263), .B2(n918), .C1(n280), .C2(n919), .A(n1050), 
        .ZN(n1045) );
  AOI22_X1 U1395 ( .A1(n921), .A2(\regOut[27][3] ), .B1(n922), .B2(
        \regOut[26][3] ), .ZN(n1050) );
  INV_X1 U1396 ( .A(\regOut[24][3] ), .ZN(n280) );
  INV_X1 U1397 ( .A(\regOut[25][3] ), .ZN(n263) );
  OAI221_X1 U1398 ( .B1(n144), .B2(n923), .C1(n161), .C2(n924), .A(n1051), 
        .ZN(n1044) );
  AOI22_X1 U1399 ( .A1(n926), .A2(\regOut[29][3] ), .B1(n927), .B2(
        \regOut[28][3] ), .ZN(n1051) );
  INV_X1 U1400 ( .A(\regOut[30][3] ), .ZN(n161) );
  INV_X1 U1401 ( .A(\regOut[31][3] ), .ZN(n144) );
  NOR4_X1 U1402 ( .A1(n1052), .A2(n1053), .A3(n1054), .A4(n1055), .ZN(n1042)
         );
  OAI221_X1 U1403 ( .B1(n365), .B2(n932), .C1(n552), .C2(n933), .A(n1056), 
        .ZN(n1055) );
  AOI22_X1 U1404 ( .A1(n935), .A2(\regOut[3][3] ), .B1(n936), .B2(
        \regOut[2][3] ), .ZN(n1056) );
  INV_X1 U1405 ( .A(\regOut[0][3] ), .ZN(n552) );
  INV_X1 U1406 ( .A(\regOut[1][3] ), .ZN(n365) );
  OAI221_X1 U1407 ( .B1(n93), .B2(n937), .C1(n110), .C2(n938), .A(n1057), .ZN(
        n1054) );
  AOI22_X1 U1408 ( .A1(n940), .A2(\regOut[7][3] ), .B1(n941), .B2(
        \regOut[6][3] ), .ZN(n1057) );
  INV_X1 U1409 ( .A(\regOut[4][3] ), .ZN(n110) );
  INV_X1 U1410 ( .A(\regOut[5][3] ), .ZN(n93) );
  OAI221_X1 U1411 ( .B1(n16), .B2(n942), .C1(n42), .C2(n943), .A(n1058), .ZN(
        n1053) );
  AOI22_X1 U1412 ( .A1(n945), .A2(\regOut[11][3] ), .B1(n946), .B2(
        \regOut[10][3] ), .ZN(n1058) );
  INV_X1 U1413 ( .A(\regOut[8][3] ), .ZN(n42) );
  INV_X1 U1414 ( .A(\regOut[9][3] ), .ZN(n16) );
  OAI221_X1 U1415 ( .B1(n484), .B2(n947), .C1(n501), .C2(n948), .A(n1059), 
        .ZN(n1052) );
  AOI22_X1 U1416 ( .A1(n950), .A2(\regOut[15][3] ), .B1(n951), .B2(
        \regOut[14][3] ), .ZN(n1059) );
  INV_X1 U1417 ( .A(\regOut[12][3] ), .ZN(n501) );
  INV_X1 U1418 ( .A(\regOut[13][3] ), .ZN(n484) );
  NAND2_X1 U1419 ( .A1(n1060), .A2(n1061), .ZN(outA[2]) );
  NOR4_X1 U1420 ( .A1(n1062), .A2(n1063), .A3(n1064), .A4(n1065), .ZN(n1061)
         );
  OAI221_X1 U1421 ( .B1(n417), .B2(n908), .C1(n434), .C2(n909), .A(n1066), 
        .ZN(n1065) );
  AOI22_X1 U1422 ( .A1(n911), .A2(\regOut[19][2] ), .B1(n912), .B2(
        \regOut[18][2] ), .ZN(n1066) );
  INV_X1 U1423 ( .A(\regOut[16][2] ), .ZN(n434) );
  INV_X1 U1424 ( .A(\regOut[17][2] ), .ZN(n417) );
  OAI221_X1 U1425 ( .B1(n332), .B2(n913), .C1(n349), .C2(n914), .A(n1067), 
        .ZN(n1064) );
  AOI22_X1 U1426 ( .A1(n916), .A2(\regOut[23][2] ), .B1(n917), .B2(
        \regOut[22][2] ), .ZN(n1067) );
  INV_X1 U1427 ( .A(\regOut[20][2] ), .ZN(n349) );
  INV_X1 U1428 ( .A(\regOut[21][2] ), .ZN(n332) );
  OAI221_X1 U1429 ( .B1(n264), .B2(n918), .C1(n281), .C2(n919), .A(n1068), 
        .ZN(n1063) );
  AOI22_X1 U1430 ( .A1(n921), .A2(\regOut[27][2] ), .B1(n922), .B2(
        \regOut[26][2] ), .ZN(n1068) );
  INV_X1 U1431 ( .A(\regOut[24][2] ), .ZN(n281) );
  INV_X1 U1432 ( .A(\regOut[25][2] ), .ZN(n264) );
  OAI221_X1 U1433 ( .B1(n145), .B2(n923), .C1(n162), .C2(n924), .A(n1069), 
        .ZN(n1062) );
  AOI22_X1 U1434 ( .A1(n926), .A2(\regOut[29][2] ), .B1(n927), .B2(
        \regOut[28][2] ), .ZN(n1069) );
  INV_X1 U1435 ( .A(\regOut[30][2] ), .ZN(n162) );
  INV_X1 U1436 ( .A(\regOut[31][2] ), .ZN(n145) );
  NOR4_X1 U1437 ( .A1(n1070), .A2(n1071), .A3(n1072), .A4(n1073), .ZN(n1060)
         );
  OAI221_X1 U1438 ( .B1(n366), .B2(n932), .C1(n553), .C2(n933), .A(n1074), 
        .ZN(n1073) );
  AOI22_X1 U1439 ( .A1(n935), .A2(\regOut[3][2] ), .B1(n936), .B2(
        \regOut[2][2] ), .ZN(n1074) );
  INV_X1 U1440 ( .A(\regOut[0][2] ), .ZN(n553) );
  INV_X1 U1441 ( .A(\regOut[1][2] ), .ZN(n366) );
  OAI221_X1 U1442 ( .B1(n94), .B2(n937), .C1(n111), .C2(n938), .A(n1075), .ZN(
        n1072) );
  AOI22_X1 U1443 ( .A1(n940), .A2(\regOut[7][2] ), .B1(n941), .B2(
        \regOut[6][2] ), .ZN(n1075) );
  INV_X1 U1444 ( .A(\regOut[4][2] ), .ZN(n111) );
  INV_X1 U1445 ( .A(\regOut[5][2] ), .ZN(n94) );
  OAI221_X1 U1446 ( .B1(n18), .B2(n942), .C1(n43), .C2(n943), .A(n1076), .ZN(
        n1071) );
  AOI22_X1 U1447 ( .A1(n945), .A2(\regOut[11][2] ), .B1(n946), .B2(
        \regOut[10][2] ), .ZN(n1076) );
  INV_X1 U1448 ( .A(\regOut[8][2] ), .ZN(n43) );
  INV_X1 U1449 ( .A(\regOut[9][2] ), .ZN(n18) );
  OAI221_X1 U1450 ( .B1(n485), .B2(n947), .C1(n502), .C2(n948), .A(n1077), 
        .ZN(n1070) );
  AOI22_X1 U1451 ( .A1(n950), .A2(\regOut[15][2] ), .B1(n951), .B2(
        \regOut[14][2] ), .ZN(n1077) );
  INV_X1 U1452 ( .A(\regOut[12][2] ), .ZN(n502) );
  INV_X1 U1453 ( .A(\regOut[13][2] ), .ZN(n485) );
  NAND2_X1 U1454 ( .A1(n1078), .A2(n1079), .ZN(outA[1]) );
  NOR4_X1 U1455 ( .A1(n1080), .A2(n1081), .A3(n1082), .A4(n1083), .ZN(n1079)
         );
  OAI221_X1 U1456 ( .B1(n418), .B2(n908), .C1(n435), .C2(n909), .A(n1084), 
        .ZN(n1083) );
  AOI22_X1 U1457 ( .A1(n911), .A2(\regOut[19][1] ), .B1(n912), .B2(
        \regOut[18][1] ), .ZN(n1084) );
  INV_X1 U1458 ( .A(\regOut[16][1] ), .ZN(n435) );
  INV_X1 U1459 ( .A(\regOut[17][1] ), .ZN(n418) );
  OAI221_X1 U1460 ( .B1(n333), .B2(n913), .C1(n350), .C2(n914), .A(n1085), 
        .ZN(n1082) );
  AOI22_X1 U1461 ( .A1(n916), .A2(\regOut[23][1] ), .B1(n917), .B2(
        \regOut[22][1] ), .ZN(n1085) );
  INV_X1 U1462 ( .A(\regOut[20][1] ), .ZN(n350) );
  INV_X1 U1463 ( .A(\regOut[21][1] ), .ZN(n333) );
  OAI221_X1 U1464 ( .B1(n265), .B2(n918), .C1(n282), .C2(n919), .A(n1086), 
        .ZN(n1081) );
  AOI22_X1 U1465 ( .A1(n921), .A2(\regOut[27][1] ), .B1(n922), .B2(
        \regOut[26][1] ), .ZN(n1086) );
  INV_X1 U1466 ( .A(\regOut[24][1] ), .ZN(n282) );
  INV_X1 U1467 ( .A(\regOut[25][1] ), .ZN(n265) );
  OAI221_X1 U1468 ( .B1(n146), .B2(n923), .C1(n163), .C2(n924), .A(n1087), 
        .ZN(n1080) );
  AOI22_X1 U1469 ( .A1(n926), .A2(\regOut[29][1] ), .B1(n927), .B2(
        \regOut[28][1] ), .ZN(n1087) );
  INV_X1 U1470 ( .A(\regOut[30][1] ), .ZN(n163) );
  INV_X1 U1471 ( .A(\regOut[31][1] ), .ZN(n146) );
  NOR4_X1 U1472 ( .A1(n1088), .A2(n1089), .A3(n1090), .A4(n1091), .ZN(n1078)
         );
  OAI221_X1 U1473 ( .B1(n367), .B2(n932), .C1(n554), .C2(n933), .A(n1092), 
        .ZN(n1091) );
  AOI22_X1 U1474 ( .A1(n935), .A2(\regOut[3][1] ), .B1(n936), .B2(
        \regOut[2][1] ), .ZN(n1092) );
  INV_X1 U1475 ( .A(\regOut[0][1] ), .ZN(n554) );
  INV_X1 U1476 ( .A(\regOut[1][1] ), .ZN(n367) );
  OAI221_X1 U1477 ( .B1(n95), .B2(n937), .C1(n112), .C2(n938), .A(n1093), .ZN(
        n1090) );
  AOI22_X1 U1478 ( .A1(n940), .A2(\regOut[7][1] ), .B1(n941), .B2(
        \regOut[6][1] ), .ZN(n1093) );
  INV_X1 U1479 ( .A(\regOut[4][1] ), .ZN(n112) );
  INV_X1 U1480 ( .A(\regOut[5][1] ), .ZN(n95) );
  OAI221_X1 U1481 ( .B1(n20), .B2(n942), .C1(n44), .C2(n943), .A(n1094), .ZN(
        n1089) );
  AOI22_X1 U1482 ( .A1(n945), .A2(\regOut[11][1] ), .B1(n946), .B2(
        \regOut[10][1] ), .ZN(n1094) );
  INV_X1 U1483 ( .A(\regOut[8][1] ), .ZN(n44) );
  INV_X1 U1484 ( .A(\regOut[9][1] ), .ZN(n20) );
  OAI221_X1 U1485 ( .B1(n486), .B2(n947), .C1(n503), .C2(n948), .A(n1095), 
        .ZN(n1088) );
  AOI22_X1 U1486 ( .A1(n950), .A2(\regOut[15][1] ), .B1(n951), .B2(
        \regOut[14][1] ), .ZN(n1095) );
  INV_X1 U1487 ( .A(\regOut[12][1] ), .ZN(n503) );
  INV_X1 U1488 ( .A(\regOut[13][1] ), .ZN(n486) );
  NAND2_X1 U1489 ( .A1(n1096), .A2(n1097), .ZN(outA[15]) );
  NOR4_X1 U1490 ( .A1(n1098), .A2(n1099), .A3(n1100), .A4(n1101), .ZN(n1097)
         );
  OAI221_X1 U1491 ( .B1(n419), .B2(n908), .C1(n436), .C2(n909), .A(n1102), 
        .ZN(n1101) );
  AOI22_X1 U1492 ( .A1(n911), .A2(\regOut[19][15] ), .B1(n912), .B2(
        \regOut[18][15] ), .ZN(n1102) );
  INV_X1 U1493 ( .A(\regOut[16][15] ), .ZN(n436) );
  INV_X1 U1494 ( .A(\regOut[17][15] ), .ZN(n419) );
  OAI221_X1 U1495 ( .B1(n334), .B2(n913), .C1(n351), .C2(n914), .A(n1103), 
        .ZN(n1100) );
  AOI22_X1 U1496 ( .A1(n916), .A2(\regOut[23][15] ), .B1(n917), .B2(
        \regOut[22][15] ), .ZN(n1103) );
  INV_X1 U1497 ( .A(\regOut[20][15] ), .ZN(n351) );
  INV_X1 U1498 ( .A(\regOut[21][15] ), .ZN(n334) );
  OAI221_X1 U1499 ( .B1(n266), .B2(n918), .C1(n283), .C2(n919), .A(n1104), 
        .ZN(n1099) );
  AOI22_X1 U1500 ( .A1(n921), .A2(\regOut[27][15] ), .B1(n922), .B2(
        \regOut[26][15] ), .ZN(n1104) );
  INV_X1 U1501 ( .A(\regOut[24][15] ), .ZN(n283) );
  INV_X1 U1502 ( .A(\regOut[25][15] ), .ZN(n266) );
  OAI221_X1 U1503 ( .B1(n147), .B2(n923), .C1(n164), .C2(n924), .A(n1105), 
        .ZN(n1098) );
  AOI22_X1 U1504 ( .A1(n926), .A2(\regOut[29][15] ), .B1(n927), .B2(
        \regOut[28][15] ), .ZN(n1105) );
  INV_X1 U1505 ( .A(\regOut[30][15] ), .ZN(n164) );
  INV_X1 U1506 ( .A(\regOut[31][15] ), .ZN(n147) );
  NOR4_X1 U1507 ( .A1(n1106), .A2(n1107), .A3(n1108), .A4(n1109), .ZN(n1096)
         );
  OAI221_X1 U1508 ( .B1(n368), .B2(n932), .C1(n555), .C2(n933), .A(n1110), 
        .ZN(n1109) );
  AOI22_X1 U1509 ( .A1(n935), .A2(\regOut[3][15] ), .B1(n936), .B2(
        \regOut[2][15] ), .ZN(n1110) );
  INV_X1 U1510 ( .A(\regOut[0][15] ), .ZN(n555) );
  INV_X1 U1511 ( .A(\regOut[1][15] ), .ZN(n368) );
  OAI221_X1 U1512 ( .B1(n96), .B2(n937), .C1(n113), .C2(n938), .A(n1111), .ZN(
        n1108) );
  AOI22_X1 U1513 ( .A1(n940), .A2(\regOut[7][15] ), .B1(n941), .B2(
        \regOut[6][15] ), .ZN(n1111) );
  INV_X1 U1514 ( .A(\regOut[4][15] ), .ZN(n113) );
  INV_X1 U1515 ( .A(\regOut[5][15] ), .ZN(n96) );
  OAI221_X1 U1516 ( .B1(n22), .B2(n942), .C1(n45), .C2(n943), .A(n1112), .ZN(
        n1107) );
  AOI22_X1 U1517 ( .A1(n945), .A2(\regOut[11][15] ), .B1(n946), .B2(
        \regOut[10][15] ), .ZN(n1112) );
  INV_X1 U1518 ( .A(\regOut[8][15] ), .ZN(n45) );
  INV_X1 U1519 ( .A(\regOut[9][15] ), .ZN(n22) );
  OAI221_X1 U1520 ( .B1(n487), .B2(n947), .C1(n504), .C2(n948), .A(n1113), 
        .ZN(n1106) );
  AOI22_X1 U1521 ( .A1(n950), .A2(\regOut[15][15] ), .B1(n951), .B2(
        \regOut[14][15] ), .ZN(n1113) );
  INV_X1 U1522 ( .A(\regOut[12][15] ), .ZN(n504) );
  INV_X1 U1523 ( .A(\regOut[13][15] ), .ZN(n487) );
  NAND2_X1 U1524 ( .A1(n1114), .A2(n1115), .ZN(outA[14]) );
  NOR4_X1 U1525 ( .A1(n1116), .A2(n1117), .A3(n1118), .A4(n1119), .ZN(n1115)
         );
  OAI221_X1 U1526 ( .B1(n420), .B2(n908), .C1(n437), .C2(n909), .A(n1120), 
        .ZN(n1119) );
  AOI22_X1 U1527 ( .A1(n911), .A2(\regOut[19][14] ), .B1(n912), .B2(
        \regOut[18][14] ), .ZN(n1120) );
  INV_X1 U1528 ( .A(\regOut[16][14] ), .ZN(n437) );
  INV_X1 U1529 ( .A(\regOut[17][14] ), .ZN(n420) );
  OAI221_X1 U1530 ( .B1(n335), .B2(n913), .C1(n352), .C2(n914), .A(n1121), 
        .ZN(n1118) );
  AOI22_X1 U1531 ( .A1(n916), .A2(\regOut[23][14] ), .B1(n917), .B2(
        \regOut[22][14] ), .ZN(n1121) );
  INV_X1 U1532 ( .A(\regOut[20][14] ), .ZN(n352) );
  INV_X1 U1533 ( .A(\regOut[21][14] ), .ZN(n335) );
  OAI221_X1 U1534 ( .B1(n267), .B2(n918), .C1(n284), .C2(n919), .A(n1122), 
        .ZN(n1117) );
  AOI22_X1 U1535 ( .A1(n921), .A2(\regOut[27][14] ), .B1(n922), .B2(
        \regOut[26][14] ), .ZN(n1122) );
  INV_X1 U1536 ( .A(\regOut[24][14] ), .ZN(n284) );
  INV_X1 U1537 ( .A(\regOut[25][14] ), .ZN(n267) );
  OAI221_X1 U1538 ( .B1(n148), .B2(n923), .C1(n165), .C2(n924), .A(n1123), 
        .ZN(n1116) );
  AOI22_X1 U1539 ( .A1(n926), .A2(\regOut[29][14] ), .B1(n927), .B2(
        \regOut[28][14] ), .ZN(n1123) );
  INV_X1 U1540 ( .A(\regOut[30][14] ), .ZN(n165) );
  INV_X1 U1541 ( .A(\regOut[31][14] ), .ZN(n148) );
  NOR4_X1 U1542 ( .A1(n1124), .A2(n1125), .A3(n1126), .A4(n1127), .ZN(n1114)
         );
  OAI221_X1 U1543 ( .B1(n369), .B2(n932), .C1(n556), .C2(n933), .A(n1128), 
        .ZN(n1127) );
  AOI22_X1 U1544 ( .A1(n935), .A2(\regOut[3][14] ), .B1(n936), .B2(
        \regOut[2][14] ), .ZN(n1128) );
  INV_X1 U1545 ( .A(\regOut[0][14] ), .ZN(n556) );
  INV_X1 U1546 ( .A(\regOut[1][14] ), .ZN(n369) );
  OAI221_X1 U1547 ( .B1(n97), .B2(n937), .C1(n114), .C2(n938), .A(n1129), .ZN(
        n1126) );
  AOI22_X1 U1548 ( .A1(n940), .A2(\regOut[7][14] ), .B1(n941), .B2(
        \regOut[6][14] ), .ZN(n1129) );
  INV_X1 U1549 ( .A(\regOut[4][14] ), .ZN(n114) );
  INV_X1 U1550 ( .A(\regOut[5][14] ), .ZN(n97) );
  OAI221_X1 U1551 ( .B1(n24), .B2(n942), .C1(n46), .C2(n943), .A(n1130), .ZN(
        n1125) );
  AOI22_X1 U1552 ( .A1(n945), .A2(\regOut[11][14] ), .B1(n946), .B2(
        \regOut[10][14] ), .ZN(n1130) );
  INV_X1 U1553 ( .A(\regOut[8][14] ), .ZN(n46) );
  INV_X1 U1554 ( .A(\regOut[9][14] ), .ZN(n24) );
  OAI221_X1 U1555 ( .B1(n488), .B2(n947), .C1(n505), .C2(n948), .A(n1131), 
        .ZN(n1124) );
  AOI22_X1 U1556 ( .A1(n950), .A2(\regOut[15][14] ), .B1(n951), .B2(
        \regOut[14][14] ), .ZN(n1131) );
  INV_X1 U1557 ( .A(\regOut[12][14] ), .ZN(n505) );
  INV_X1 U1558 ( .A(\regOut[13][14] ), .ZN(n488) );
  NAND2_X1 U1559 ( .A1(n1132), .A2(n1133), .ZN(outA[13]) );
  NOR4_X1 U1560 ( .A1(n1134), .A2(n1135), .A3(n1136), .A4(n1137), .ZN(n1133)
         );
  OAI221_X1 U1561 ( .B1(n421), .B2(n908), .C1(n438), .C2(n909), .A(n1138), 
        .ZN(n1137) );
  AOI22_X1 U1562 ( .A1(n911), .A2(\regOut[19][13] ), .B1(n912), .B2(
        \regOut[18][13] ), .ZN(n1138) );
  INV_X1 U1563 ( .A(\regOut[16][13] ), .ZN(n438) );
  INV_X1 U1564 ( .A(\regOut[17][13] ), .ZN(n421) );
  OAI221_X1 U1565 ( .B1(n336), .B2(n913), .C1(n353), .C2(n914), .A(n1139), 
        .ZN(n1136) );
  AOI22_X1 U1566 ( .A1(n916), .A2(\regOut[23][13] ), .B1(n917), .B2(
        \regOut[22][13] ), .ZN(n1139) );
  INV_X1 U1567 ( .A(\regOut[20][13] ), .ZN(n353) );
  INV_X1 U1568 ( .A(\regOut[21][13] ), .ZN(n336) );
  OAI221_X1 U1569 ( .B1(n268), .B2(n918), .C1(n285), .C2(n919), .A(n1140), 
        .ZN(n1135) );
  AOI22_X1 U1570 ( .A1(n921), .A2(\regOut[27][13] ), .B1(n922), .B2(
        \regOut[26][13] ), .ZN(n1140) );
  INV_X1 U1571 ( .A(\regOut[24][13] ), .ZN(n285) );
  INV_X1 U1572 ( .A(\regOut[25][13] ), .ZN(n268) );
  OAI221_X1 U1573 ( .B1(n149), .B2(n923), .C1(n166), .C2(n924), .A(n1141), 
        .ZN(n1134) );
  AOI22_X1 U1574 ( .A1(n926), .A2(\regOut[29][13] ), .B1(n927), .B2(
        \regOut[28][13] ), .ZN(n1141) );
  INV_X1 U1575 ( .A(\regOut[30][13] ), .ZN(n166) );
  INV_X1 U1576 ( .A(\regOut[31][13] ), .ZN(n149) );
  NOR4_X1 U1577 ( .A1(n1142), .A2(n1143), .A3(n1144), .A4(n1145), .ZN(n1132)
         );
  OAI221_X1 U1578 ( .B1(n370), .B2(n932), .C1(n557), .C2(n933), .A(n1146), 
        .ZN(n1145) );
  AOI22_X1 U1579 ( .A1(n935), .A2(\regOut[3][13] ), .B1(n936), .B2(
        \regOut[2][13] ), .ZN(n1146) );
  INV_X1 U1580 ( .A(\regOut[0][13] ), .ZN(n557) );
  INV_X1 U1581 ( .A(\regOut[1][13] ), .ZN(n370) );
  OAI221_X1 U1582 ( .B1(n98), .B2(n937), .C1(n115), .C2(n938), .A(n1147), .ZN(
        n1144) );
  AOI22_X1 U1583 ( .A1(n940), .A2(\regOut[7][13] ), .B1(n941), .B2(
        \regOut[6][13] ), .ZN(n1147) );
  INV_X1 U1584 ( .A(\regOut[4][13] ), .ZN(n115) );
  INV_X1 U1585 ( .A(\regOut[5][13] ), .ZN(n98) );
  OAI221_X1 U1586 ( .B1(n26), .B2(n942), .C1(n47), .C2(n943), .A(n1148), .ZN(
        n1143) );
  AOI22_X1 U1587 ( .A1(n945), .A2(\regOut[11][13] ), .B1(n946), .B2(
        \regOut[10][13] ), .ZN(n1148) );
  INV_X1 U1588 ( .A(\regOut[8][13] ), .ZN(n47) );
  INV_X1 U1589 ( .A(\regOut[9][13] ), .ZN(n26) );
  OAI221_X1 U1590 ( .B1(n489), .B2(n947), .C1(n506), .C2(n948), .A(n1149), 
        .ZN(n1142) );
  AOI22_X1 U1591 ( .A1(n950), .A2(\regOut[15][13] ), .B1(n951), .B2(
        \regOut[14][13] ), .ZN(n1149) );
  INV_X1 U1592 ( .A(\regOut[12][13] ), .ZN(n506) );
  INV_X1 U1593 ( .A(\regOut[13][13] ), .ZN(n489) );
  NAND2_X1 U1594 ( .A1(n1150), .A2(n1151), .ZN(outA[12]) );
  NOR4_X1 U1595 ( .A1(n1152), .A2(n1153), .A3(n1154), .A4(n1155), .ZN(n1151)
         );
  OAI221_X1 U1596 ( .B1(n422), .B2(n908), .C1(n439), .C2(n909), .A(n1156), 
        .ZN(n1155) );
  AOI22_X1 U1597 ( .A1(n911), .A2(\regOut[19][12] ), .B1(n912), .B2(
        \regOut[18][12] ), .ZN(n1156) );
  INV_X1 U1598 ( .A(\regOut[16][12] ), .ZN(n439) );
  INV_X1 U1599 ( .A(\regOut[17][12] ), .ZN(n422) );
  OAI221_X1 U1600 ( .B1(n337), .B2(n913), .C1(n354), .C2(n914), .A(n1157), 
        .ZN(n1154) );
  AOI22_X1 U1601 ( .A1(n916), .A2(\regOut[23][12] ), .B1(n917), .B2(
        \regOut[22][12] ), .ZN(n1157) );
  INV_X1 U1602 ( .A(\regOut[20][12] ), .ZN(n354) );
  INV_X1 U1603 ( .A(\regOut[21][12] ), .ZN(n337) );
  OAI221_X1 U1604 ( .B1(n269), .B2(n918), .C1(n286), .C2(n919), .A(n1158), 
        .ZN(n1153) );
  AOI22_X1 U1605 ( .A1(n921), .A2(\regOut[27][12] ), .B1(n922), .B2(
        \regOut[26][12] ), .ZN(n1158) );
  INV_X1 U1606 ( .A(\regOut[24][12] ), .ZN(n286) );
  INV_X1 U1607 ( .A(\regOut[25][12] ), .ZN(n269) );
  OAI221_X1 U1608 ( .B1(n150), .B2(n923), .C1(n167), .C2(n924), .A(n1159), 
        .ZN(n1152) );
  AOI22_X1 U1609 ( .A1(n926), .A2(\regOut[29][12] ), .B1(n927), .B2(
        \regOut[28][12] ), .ZN(n1159) );
  INV_X1 U1610 ( .A(\regOut[30][12] ), .ZN(n167) );
  INV_X1 U1611 ( .A(\regOut[31][12] ), .ZN(n150) );
  NOR4_X1 U1612 ( .A1(n1160), .A2(n1161), .A3(n1162), .A4(n1163), .ZN(n1150)
         );
  OAI221_X1 U1613 ( .B1(n371), .B2(n932), .C1(n558), .C2(n933), .A(n1164), 
        .ZN(n1163) );
  AOI22_X1 U1614 ( .A1(n935), .A2(\regOut[3][12] ), .B1(n936), .B2(
        \regOut[2][12] ), .ZN(n1164) );
  INV_X1 U1615 ( .A(\regOut[0][12] ), .ZN(n558) );
  INV_X1 U1616 ( .A(\regOut[1][12] ), .ZN(n371) );
  OAI221_X1 U1617 ( .B1(n99), .B2(n937), .C1(n116), .C2(n938), .A(n1165), .ZN(
        n1162) );
  AOI22_X1 U1618 ( .A1(n940), .A2(\regOut[7][12] ), .B1(n941), .B2(
        \regOut[6][12] ), .ZN(n1165) );
  INV_X1 U1619 ( .A(\regOut[4][12] ), .ZN(n116) );
  INV_X1 U1620 ( .A(\regOut[5][12] ), .ZN(n99) );
  OAI221_X1 U1621 ( .B1(n28), .B2(n942), .C1(n48), .C2(n943), .A(n1166), .ZN(
        n1161) );
  AOI22_X1 U1622 ( .A1(n945), .A2(\regOut[11][12] ), .B1(n946), .B2(
        \regOut[10][12] ), .ZN(n1166) );
  INV_X1 U1623 ( .A(\regOut[8][12] ), .ZN(n48) );
  INV_X1 U1624 ( .A(\regOut[9][12] ), .ZN(n28) );
  OAI221_X1 U1625 ( .B1(n490), .B2(n947), .C1(n507), .C2(n948), .A(n1167), 
        .ZN(n1160) );
  AOI22_X1 U1626 ( .A1(n950), .A2(\regOut[15][12] ), .B1(n951), .B2(
        \regOut[14][12] ), .ZN(n1167) );
  INV_X1 U1627 ( .A(\regOut[12][12] ), .ZN(n507) );
  INV_X1 U1628 ( .A(\regOut[13][12] ), .ZN(n490) );
  NAND2_X1 U1629 ( .A1(n1168), .A2(n1169), .ZN(outA[11]) );
  NOR4_X1 U1630 ( .A1(n1170), .A2(n1171), .A3(n1172), .A4(n1173), .ZN(n1169)
         );
  OAI221_X1 U1631 ( .B1(n423), .B2(n908), .C1(n440), .C2(n909), .A(n1174), 
        .ZN(n1173) );
  AOI22_X1 U1632 ( .A1(n911), .A2(\regOut[19][11] ), .B1(n912), .B2(
        \regOut[18][11] ), .ZN(n1174) );
  INV_X1 U1633 ( .A(\regOut[16][11] ), .ZN(n440) );
  INV_X1 U1634 ( .A(\regOut[17][11] ), .ZN(n423) );
  OAI221_X1 U1635 ( .B1(n338), .B2(n913), .C1(n355), .C2(n914), .A(n1175), 
        .ZN(n1172) );
  AOI22_X1 U1636 ( .A1(n916), .A2(\regOut[23][11] ), .B1(n917), .B2(
        \regOut[22][11] ), .ZN(n1175) );
  INV_X1 U1637 ( .A(\regOut[20][11] ), .ZN(n355) );
  INV_X1 U1638 ( .A(\regOut[21][11] ), .ZN(n338) );
  OAI221_X1 U1639 ( .B1(n270), .B2(n918), .C1(n287), .C2(n919), .A(n1176), 
        .ZN(n1171) );
  AOI22_X1 U1640 ( .A1(n921), .A2(\regOut[27][11] ), .B1(n922), .B2(
        \regOut[26][11] ), .ZN(n1176) );
  INV_X1 U1641 ( .A(\regOut[24][11] ), .ZN(n287) );
  INV_X1 U1642 ( .A(\regOut[25][11] ), .ZN(n270) );
  OAI221_X1 U1643 ( .B1(n151), .B2(n923), .C1(n168), .C2(n924), .A(n1177), 
        .ZN(n1170) );
  AOI22_X1 U1644 ( .A1(n926), .A2(\regOut[29][11] ), .B1(n927), .B2(
        \regOut[28][11] ), .ZN(n1177) );
  INV_X1 U1645 ( .A(\regOut[30][11] ), .ZN(n168) );
  INV_X1 U1646 ( .A(\regOut[31][11] ), .ZN(n151) );
  NOR4_X1 U1647 ( .A1(n1178), .A2(n1179), .A3(n1180), .A4(n1181), .ZN(n1168)
         );
  OAI221_X1 U1648 ( .B1(n372), .B2(n932), .C1(n559), .C2(n933), .A(n1182), 
        .ZN(n1181) );
  AOI22_X1 U1649 ( .A1(n935), .A2(\regOut[3][11] ), .B1(n936), .B2(
        \regOut[2][11] ), .ZN(n1182) );
  INV_X1 U1650 ( .A(\regOut[0][11] ), .ZN(n559) );
  INV_X1 U1651 ( .A(\regOut[1][11] ), .ZN(n372) );
  OAI221_X1 U1652 ( .B1(n100), .B2(n937), .C1(n117), .C2(n938), .A(n1183), 
        .ZN(n1180) );
  AOI22_X1 U1653 ( .A1(n940), .A2(\regOut[7][11] ), .B1(n941), .B2(
        \regOut[6][11] ), .ZN(n1183) );
  INV_X1 U1654 ( .A(\regOut[4][11] ), .ZN(n117) );
  INV_X1 U1655 ( .A(\regOut[5][11] ), .ZN(n100) );
  OAI221_X1 U1656 ( .B1(n30), .B2(n942), .C1(n49), .C2(n943), .A(n1184), .ZN(
        n1179) );
  AOI22_X1 U1657 ( .A1(n945), .A2(\regOut[11][11] ), .B1(n946), .B2(
        \regOut[10][11] ), .ZN(n1184) );
  INV_X1 U1658 ( .A(\regOut[8][11] ), .ZN(n49) );
  INV_X1 U1659 ( .A(\regOut[9][11] ), .ZN(n30) );
  OAI221_X1 U1660 ( .B1(n491), .B2(n947), .C1(n508), .C2(n948), .A(n1185), 
        .ZN(n1178) );
  AOI22_X1 U1661 ( .A1(n950), .A2(\regOut[15][11] ), .B1(n951), .B2(
        \regOut[14][11] ), .ZN(n1185) );
  INV_X1 U1662 ( .A(\regOut[12][11] ), .ZN(n508) );
  INV_X1 U1663 ( .A(\regOut[13][11] ), .ZN(n491) );
  NAND2_X1 U1664 ( .A1(n1186), .A2(n1187), .ZN(outA[10]) );
  NOR4_X1 U1665 ( .A1(n1188), .A2(n1189), .A3(n1190), .A4(n1191), .ZN(n1187)
         );
  OAI221_X1 U1666 ( .B1(n424), .B2(n908), .C1(n441), .C2(n909), .A(n1192), 
        .ZN(n1191) );
  AOI22_X1 U1667 ( .A1(n911), .A2(\regOut[19][10] ), .B1(n912), .B2(
        \regOut[18][10] ), .ZN(n1192) );
  INV_X1 U1668 ( .A(\regOut[16][10] ), .ZN(n441) );
  INV_X1 U1669 ( .A(\regOut[17][10] ), .ZN(n424) );
  OAI221_X1 U1670 ( .B1(n339), .B2(n913), .C1(n356), .C2(n914), .A(n1193), 
        .ZN(n1190) );
  AOI22_X1 U1671 ( .A1(n916), .A2(\regOut[23][10] ), .B1(n917), .B2(
        \regOut[22][10] ), .ZN(n1193) );
  INV_X1 U1672 ( .A(\regOut[20][10] ), .ZN(n356) );
  INV_X1 U1673 ( .A(\regOut[21][10] ), .ZN(n339) );
  OAI221_X1 U1674 ( .B1(n271), .B2(n918), .C1(n288), .C2(n919), .A(n1194), 
        .ZN(n1189) );
  AOI22_X1 U1675 ( .A1(n921), .A2(\regOut[27][10] ), .B1(n922), .B2(
        \regOut[26][10] ), .ZN(n1194) );
  INV_X1 U1676 ( .A(\regOut[24][10] ), .ZN(n288) );
  INV_X1 U1677 ( .A(\regOut[25][10] ), .ZN(n271) );
  OAI221_X1 U1678 ( .B1(n152), .B2(n923), .C1(n169), .C2(n924), .A(n1195), 
        .ZN(n1188) );
  AOI22_X1 U1679 ( .A1(n926), .A2(\regOut[29][10] ), .B1(n927), .B2(
        \regOut[28][10] ), .ZN(n1195) );
  INV_X1 U1680 ( .A(\regOut[30][10] ), .ZN(n169) );
  INV_X1 U1681 ( .A(\regOut[31][10] ), .ZN(n152) );
  NOR4_X1 U1682 ( .A1(n1196), .A2(n1197), .A3(n1198), .A4(n1199), .ZN(n1186)
         );
  OAI221_X1 U1683 ( .B1(n373), .B2(n932), .C1(n560), .C2(n933), .A(n1200), 
        .ZN(n1199) );
  AOI22_X1 U1684 ( .A1(n935), .A2(\regOut[3][10] ), .B1(n936), .B2(
        \regOut[2][10] ), .ZN(n1200) );
  INV_X1 U1685 ( .A(\regOut[0][10] ), .ZN(n560) );
  INV_X1 U1686 ( .A(\regOut[1][10] ), .ZN(n373) );
  OAI221_X1 U1687 ( .B1(n101), .B2(n937), .C1(n118), .C2(n938), .A(n1201), 
        .ZN(n1198) );
  AOI22_X1 U1688 ( .A1(n940), .A2(\regOut[7][10] ), .B1(n941), .B2(
        \regOut[6][10] ), .ZN(n1201) );
  INV_X1 U1689 ( .A(\regOut[4][10] ), .ZN(n118) );
  INV_X1 U1690 ( .A(\regOut[5][10] ), .ZN(n101) );
  OAI221_X1 U1691 ( .B1(n32), .B2(n942), .C1(n50), .C2(n943), .A(n1202), .ZN(
        n1197) );
  AOI22_X1 U1692 ( .A1(n945), .A2(\regOut[11][10] ), .B1(n946), .B2(
        \regOut[10][10] ), .ZN(n1202) );
  INV_X1 U1693 ( .A(\regOut[8][10] ), .ZN(n50) );
  INV_X1 U1694 ( .A(\regOut[9][10] ), .ZN(n32) );
  OAI221_X1 U1695 ( .B1(n492), .B2(n947), .C1(n509), .C2(n948), .A(n1203), 
        .ZN(n1196) );
  AOI22_X1 U1696 ( .A1(n950), .A2(\regOut[15][10] ), .B1(n951), .B2(
        \regOut[14][10] ), .ZN(n1203) );
  INV_X1 U1697 ( .A(\regOut[12][10] ), .ZN(n509) );
  INV_X1 U1698 ( .A(\regOut[13][10] ), .ZN(n492) );
  NAND2_X1 U1699 ( .A1(n1204), .A2(n1205), .ZN(outA[0]) );
  NOR4_X1 U1700 ( .A1(n1206), .A2(n1207), .A3(n1208), .A4(n1209), .ZN(n1205)
         );
  OAI221_X1 U1701 ( .B1(n425), .B2(n908), .C1(n442), .C2(n909), .A(n1210), 
        .ZN(n1209) );
  AOI22_X1 U1702 ( .A1(n911), .A2(\regOut[19][0] ), .B1(n912), .B2(
        \regOut[18][0] ), .ZN(n1210) );
  AND2_X1 U1703 ( .A1(n1211), .A2(n1212), .ZN(n912) );
  AND2_X1 U1704 ( .A1(n1213), .A2(n1212), .ZN(n911) );
  NAND2_X1 U1705 ( .A1(n1211), .A2(n1214), .ZN(n909) );
  INV_X1 U1706 ( .A(\regOut[16][0] ), .ZN(n442) );
  NAND2_X1 U1707 ( .A1(n1213), .A2(n1214), .ZN(n908) );
  INV_X1 U1708 ( .A(\regOut[17][0] ), .ZN(n425) );
  OAI221_X1 U1709 ( .B1(n340), .B2(n913), .C1(n357), .C2(n914), .A(n1215), 
        .ZN(n1208) );
  AOI22_X1 U1710 ( .A1(n916), .A2(\regOut[23][0] ), .B1(n917), .B2(
        \regOut[22][0] ), .ZN(n1215) );
  AND2_X1 U1711 ( .A1(n1211), .A2(n1216), .ZN(n917) );
  AND2_X1 U1712 ( .A1(n1213), .A2(n1216), .ZN(n916) );
  NAND2_X1 U1713 ( .A1(n1211), .A2(n1217), .ZN(n914) );
  AND2_X1 U1714 ( .A1(n1218), .A2(n1219), .ZN(n1211) );
  INV_X1 U1715 ( .A(\regOut[20][0] ), .ZN(n357) );
  NAND2_X1 U1716 ( .A1(n1213), .A2(n1217), .ZN(n913) );
  AND2_X1 U1717 ( .A1(n1218), .A2(n1250), .ZN(n1213) );
  AND2_X1 U1718 ( .A1(n1248), .A2(n1220), .ZN(n1218) );
  INV_X1 U1719 ( .A(\regOut[21][0] ), .ZN(n340) );
  OAI221_X1 U1720 ( .B1(n272), .B2(n918), .C1(n289), .C2(n919), .A(n1221), 
        .ZN(n1207) );
  AOI22_X1 U1721 ( .A1(n921), .A2(\regOut[27][0] ), .B1(n922), .B2(
        \regOut[26][0] ), .ZN(n1221) );
  AND2_X1 U1722 ( .A1(n1212), .A2(n1222), .ZN(n922) );
  AND2_X1 U1723 ( .A1(n1212), .A2(n1223), .ZN(n921) );
  NAND2_X1 U1724 ( .A1(n1214), .A2(n1222), .ZN(n919) );
  INV_X1 U1725 ( .A(\regOut[24][0] ), .ZN(n289) );
  NAND2_X1 U1726 ( .A1(n1214), .A2(n1223), .ZN(n918) );
  INV_X1 U1727 ( .A(\regOut[25][0] ), .ZN(n272) );
  OAI221_X1 U1728 ( .B1(n153), .B2(n923), .C1(n170), .C2(n924), .A(n1224), 
        .ZN(n1206) );
  AOI22_X1 U1729 ( .A1(n926), .A2(\regOut[29][0] ), .B1(n927), .B2(
        \regOut[28][0] ), .ZN(n1224) );
  AND2_X1 U1730 ( .A1(n1217), .A2(n1222), .ZN(n927) );
  AND2_X1 U1731 ( .A1(n1217), .A2(n1223), .ZN(n926) );
  NAND2_X1 U1732 ( .A1(n1222), .A2(n1216), .ZN(n924) );
  AND2_X1 U1733 ( .A1(n1225), .A2(n1219), .ZN(n1222) );
  INV_X1 U1734 ( .A(\regOut[30][0] ), .ZN(n170) );
  NAND2_X1 U1735 ( .A1(n1216), .A2(n1223), .ZN(n923) );
  AND2_X1 U1736 ( .A1(n1250), .A2(n1225), .ZN(n1223) );
  AND2_X1 U1737 ( .A1(n1248), .A2(n1246), .ZN(n1225) );
  INV_X1 U1738 ( .A(\regOut[31][0] ), .ZN(n153) );
  NOR4_X1 U1739 ( .A1(n1226), .A2(n1227), .A3(n1228), .A4(n1229), .ZN(n1204)
         );
  OAI221_X1 U1740 ( .B1(n374), .B2(n932), .C1(n561), .C2(n933), .A(n1230), 
        .ZN(n1229) );
  AOI22_X1 U1741 ( .A1(n935), .A2(\regOut[3][0] ), .B1(n936), .B2(
        \regOut[2][0] ), .ZN(n1230) );
  AND2_X1 U1742 ( .A1(n1231), .A2(n1212), .ZN(n936) );
  AND2_X1 U1743 ( .A1(n1232), .A2(n1212), .ZN(n935) );
  NAND2_X1 U1744 ( .A1(n1231), .A2(n1214), .ZN(n933) );
  INV_X1 U1745 ( .A(\regOut[0][0] ), .ZN(n561) );
  NAND2_X1 U1746 ( .A1(n1232), .A2(n1214), .ZN(n932) );
  INV_X1 U1747 ( .A(\regOut[1][0] ), .ZN(n374) );
  OAI221_X1 U1748 ( .B1(n102), .B2(n937), .C1(n119), .C2(n938), .A(n1233), 
        .ZN(n1228) );
  AOI22_X1 U1749 ( .A1(n940), .A2(\regOut[7][0] ), .B1(n941), .B2(
        \regOut[6][0] ), .ZN(n1233) );
  AND2_X1 U1750 ( .A1(n1231), .A2(n1216), .ZN(n941) );
  AND2_X1 U1751 ( .A1(n1232), .A2(n1216), .ZN(n940) );
  NAND2_X1 U1752 ( .A1(n1231), .A2(n1217), .ZN(n938) );
  AND2_X1 U1753 ( .A1(n1234), .A2(n1219), .ZN(n1231) );
  INV_X1 U1754 ( .A(\regOut[4][0] ), .ZN(n119) );
  NAND2_X1 U1755 ( .A1(n1232), .A2(n1217), .ZN(n937) );
  AND2_X1 U1756 ( .A1(n1234), .A2(n1250), .ZN(n1232) );
  NOR2_X1 U1757 ( .A1(n1246), .A2(n1248), .ZN(n1234) );
  INV_X1 U1758 ( .A(\regOut[5][0] ), .ZN(n102) );
  OAI221_X1 U1759 ( .B1(n34), .B2(n942), .C1(n51), .C2(n943), .A(n1235), .ZN(
        n1227) );
  AOI22_X1 U1760 ( .A1(n945), .A2(\regOut[11][0] ), .B1(n946), .B2(
        \regOut[10][0] ), .ZN(n1235) );
  AND2_X1 U1761 ( .A1(n1236), .A2(n1212), .ZN(n946) );
  AND2_X1 U1762 ( .A1(n1237), .A2(n1212), .ZN(n945) );
  NOR2_X1 U1763 ( .A1(n1238), .A2(n1244), .ZN(n1212) );
  NAND2_X1 U1764 ( .A1(n1236), .A2(n1214), .ZN(n943) );
  INV_X1 U1765 ( .A(\regOut[8][0] ), .ZN(n51) );
  NAND2_X1 U1766 ( .A1(n1237), .A2(n1214), .ZN(n942) );
  NOR2_X1 U1767 ( .A1(n1242), .A2(n1244), .ZN(n1214) );
  INV_X1 U1768 ( .A(\regOut[9][0] ), .ZN(n34) );
  OAI221_X1 U1769 ( .B1(n493), .B2(n947), .C1(n510), .C2(n948), .A(n1239), 
        .ZN(n1226) );
  AOI22_X1 U1770 ( .A1(n950), .A2(\regOut[15][0] ), .B1(n951), .B2(
        \regOut[14][0] ), .ZN(n1239) );
  AND2_X1 U1771 ( .A1(n1236), .A2(n1216), .ZN(n951) );
  AND2_X1 U1772 ( .A1(n1237), .A2(n1216), .ZN(n950) );
  NOR2_X1 U1773 ( .A1(n1240), .A2(n1238), .ZN(n1216) );
  INV_X1 U1774 ( .A(n1242), .ZN(n1238) );
  NAND2_X1 U1775 ( .A1(n1236), .A2(n1217), .ZN(n948) );
  AND2_X1 U1776 ( .A1(n1241), .A2(n1219), .ZN(n1236) );
  INV_X1 U1777 ( .A(n1250), .ZN(n1219) );
  INV_X1 U1778 ( .A(\regOut[12][0] ), .ZN(n510) );
  NAND2_X1 U1779 ( .A1(n1237), .A2(n1217), .ZN(n947) );
  NOR2_X1 U1780 ( .A1(n1240), .A2(n1242), .ZN(n1217) );
  INV_X1 U1781 ( .A(n1244), .ZN(n1240) );
  AND2_X1 U1782 ( .A1(n1241), .A2(n1250), .ZN(n1237) );
  NOR2_X1 U1783 ( .A1(n1220), .A2(n1248), .ZN(n1241) );
  INV_X1 U1784 ( .A(n1246), .ZN(n1220) );
  INV_X1 U1785 ( .A(\regOut[13][0] ), .ZN(n493) );
  SingleReg_31 RegX_0 ( .data({\regIn[0][15] , \regIn[0][14] , \regIn[0][13] , 
        \regIn[0][12] , \regIn[0][11] , \regIn[0][10] , \regIn[0][9] , 
        \regIn[0][8] , \regIn[0][7] , \regIn[0][6] , \regIn[0][5] , 
        \regIn[0][4] , \regIn[0][3] , \regIn[0][2] , \regIn[0][1] , 
        \regIn[0][0] }), .clk(clk), .reset(n1273), .write(n1275), .dataOut({
        \regOut[0][15] , \regOut[0][14] , \regOut[0][13] , \regOut[0][12] , 
        \regOut[0][11] , \regOut[0][10] , \regOut[0][9] , \regOut[0][8] , 
        \regOut[0][7] , \regOut[0][6] , \regOut[0][5] , \regOut[0][4] , 
        \regOut[0][3] , \regOut[0][2] , \regOut[0][1] , \regOut[0][0] }) );
  SingleReg_30 RegX_1 ( .data({\regIn[1][15] , \regIn[1][14] , \regIn[1][13] , 
        \regIn[1][12] , \regIn[1][11] , \regIn[1][10] , \regIn[1][9] , 
        \regIn[1][8] , \regIn[1][7] , \regIn[1][6] , \regIn[1][5] , 
        \regIn[1][4] , \regIn[1][3] , \regIn[1][2] , \regIn[1][1] , 
        \regIn[1][0] }), .clk(clk), .reset(n1273), .write(n1274), .dataOut({
        \regOut[1][15] , \regOut[1][14] , \regOut[1][13] , \regOut[1][12] , 
        \regOut[1][11] , \regOut[1][10] , \regOut[1][9] , \regOut[1][8] , 
        \regOut[1][7] , \regOut[1][6] , \regOut[1][5] , \regOut[1][4] , 
        \regOut[1][3] , \regOut[1][2] , \regOut[1][1] , \regOut[1][0] }) );
  SingleReg_29 RegX_2 ( .data({\regIn[2][15] , \regIn[2][14] , \regIn[2][13] , 
        \regIn[2][12] , \regIn[2][11] , \regIn[2][10] , \regIn[2][9] , 
        \regIn[2][8] , \regIn[2][7] , \regIn[2][6] , \regIn[2][5] , 
        \regIn[2][4] , \regIn[2][3] , \regIn[2][2] , \regIn[2][1] , 
        \regIn[2][0] }), .clk(clk), .reset(n1273), .write(n1274), .dataOut({
        \regOut[2][15] , \regOut[2][14] , \regOut[2][13] , \regOut[2][12] , 
        \regOut[2][11] , \regOut[2][10] , \regOut[2][9] , \regOut[2][8] , 
        \regOut[2][7] , \regOut[2][6] , \regOut[2][5] , \regOut[2][4] , 
        \regOut[2][3] , \regOut[2][2] , \regOut[2][1] , \regOut[2][0] }) );
  SingleReg_28 RegX_3 ( .data({\regIn[3][15] , \regIn[3][14] , \regIn[3][13] , 
        \regIn[3][12] , \regIn[3][11] , \regIn[3][10] , \regIn[3][9] , 
        \regIn[3][8] , \regIn[3][7] , \regIn[3][6] , \regIn[3][5] , 
        \regIn[3][4] , \regIn[3][3] , \regIn[3][2] , \regIn[3][1] , 
        \regIn[3][0] }), .clk(clk), .reset(n1273), .write(n1274), .dataOut({
        \regOut[3][15] , \regOut[3][14] , \regOut[3][13] , \regOut[3][12] , 
        \regOut[3][11] , \regOut[3][10] , \regOut[3][9] , \regOut[3][8] , 
        \regOut[3][7] , \regOut[3][6] , \regOut[3][5] , \regOut[3][4] , 
        \regOut[3][3] , \regOut[3][2] , \regOut[3][1] , \regOut[3][0] }) );
  SingleReg_27 RegX_4 ( .data({\regIn[4][15] , \regIn[4][14] , \regIn[4][13] , 
        \regIn[4][12] , \regIn[4][11] , \regIn[4][10] , \regIn[4][9] , 
        \regIn[4][8] , \regIn[4][7] , \regIn[4][6] , \regIn[4][5] , 
        \regIn[4][4] , \regIn[4][3] , \regIn[4][2] , \regIn[4][1] , 
        \regIn[4][0] }), .clk(clk), .reset(n1273), .write(n1274), .dataOut({
        \regOut[4][15] , \regOut[4][14] , \regOut[4][13] , \regOut[4][12] , 
        \regOut[4][11] , \regOut[4][10] , \regOut[4][9] , \regOut[4][8] , 
        \regOut[4][7] , \regOut[4][6] , \regOut[4][5] , \regOut[4][4] , 
        \regOut[4][3] , \regOut[4][2] , \regOut[4][1] , \regOut[4][0] }) );
  SingleReg_26 RegX_5 ( .data({\regIn[5][15] , \regIn[5][14] , \regIn[5][13] , 
        \regIn[5][12] , \regIn[5][11] , \regIn[5][10] , \regIn[5][9] , 
        \regIn[5][8] , \regIn[5][7] , \regIn[5][6] , \regIn[5][5] , 
        \regIn[5][4] , \regIn[5][3] , \regIn[5][2] , \regIn[5][1] , 
        \regIn[5][0] }), .clk(clk), .reset(n1273), .write(n1274), .dataOut({
        \regOut[5][15] , \regOut[5][14] , \regOut[5][13] , \regOut[5][12] , 
        \regOut[5][11] , \regOut[5][10] , \regOut[5][9] , \regOut[5][8] , 
        \regOut[5][7] , \regOut[5][6] , \regOut[5][5] , \regOut[5][4] , 
        \regOut[5][3] , \regOut[5][2] , \regOut[5][1] , \regOut[5][0] }) );
  SingleReg_25 RegX_6 ( .data({\regIn[6][15] , \regIn[6][14] , \regIn[6][13] , 
        \regIn[6][12] , \regIn[6][11] , \regIn[6][10] , \regIn[6][9] , 
        \regIn[6][8] , \regIn[6][7] , \regIn[6][6] , \regIn[6][5] , 
        \regIn[6][4] , \regIn[6][3] , \regIn[6][2] , \regIn[6][1] , 
        \regIn[6][0] }), .clk(clk), .reset(n1273), .write(n1274), .dataOut({
        \regOut[6][15] , \regOut[6][14] , \regOut[6][13] , \regOut[6][12] , 
        \regOut[6][11] , \regOut[6][10] , \regOut[6][9] , \regOut[6][8] , 
        \regOut[6][7] , \regOut[6][6] , \regOut[6][5] , \regOut[6][4] , 
        \regOut[6][3] , \regOut[6][2] , \regOut[6][1] , \regOut[6][0] }) );
  SingleReg_24 RegX_7 ( .data({\regIn[7][15] , \regIn[7][14] , \regIn[7][13] , 
        \regIn[7][12] , \regIn[7][11] , \regIn[7][10] , \regIn[7][9] , 
        \regIn[7][8] , \regIn[7][7] , \regIn[7][6] , \regIn[7][5] , 
        \regIn[7][4] , \regIn[7][3] , \regIn[7][2] , \regIn[7][1] , 
        \regIn[7][0] }), .clk(clk), .reset(n1273), .write(n1274), .dataOut({
        \regOut[7][15] , \regOut[7][14] , \regOut[7][13] , \regOut[7][12] , 
        \regOut[7][11] , \regOut[7][10] , \regOut[7][9] , \regOut[7][8] , 
        \regOut[7][7] , \regOut[7][6] , \regOut[7][5] , \regOut[7][4] , 
        \regOut[7][3] , \regOut[7][2] , \regOut[7][1] , \regOut[7][0] }) );
  SingleReg_23 RegX_8 ( .data({\regIn[8][15] , \regIn[8][14] , \regIn[8][13] , 
        \regIn[8][12] , \regIn[8][11] , \regIn[8][10] , \regIn[8][9] , 
        \regIn[8][8] , \regIn[8][7] , \regIn[8][6] , \regIn[8][5] , 
        \regIn[8][4] , \regIn[8][3] , \regIn[8][2] , \regIn[8][1] , 
        \regIn[8][0] }), .clk(clk), .reset(n1273), .write(n1274), .dataOut({
        \regOut[8][15] , \regOut[8][14] , \regOut[8][13] , \regOut[8][12] , 
        \regOut[8][11] , \regOut[8][10] , \regOut[8][9] , \regOut[8][8] , 
        \regOut[8][7] , \regOut[8][6] , \regOut[8][5] , \regOut[8][4] , 
        \regOut[8][3] , \regOut[8][2] , \regOut[8][1] , \regOut[8][0] }) );
  SingleReg_22 RegX_9 ( .data({\regIn[9][15] , \regIn[9][14] , \regIn[9][13] , 
        \regIn[9][12] , \regIn[9][11] , \regIn[9][10] , \regIn[9][9] , 
        \regIn[9][8] , \regIn[9][7] , \regIn[9][6] , \regIn[9][5] , 
        \regIn[9][4] , \regIn[9][3] , \regIn[9][2] , \regIn[9][1] , 
        \regIn[9][0] }), .clk(clk), .reset(n1273), .write(n1274), .dataOut({
        \regOut[9][15] , \regOut[9][14] , \regOut[9][13] , \regOut[9][12] , 
        \regOut[9][11] , \regOut[9][10] , \regOut[9][9] , \regOut[9][8] , 
        \regOut[9][7] , \regOut[9][6] , \regOut[9][5] , \regOut[9][4] , 
        \regOut[9][3] , \regOut[9][2] , \regOut[9][1] , \regOut[9][0] }) );
  SingleReg_21 RegX_10 ( .data({\regIn[10][15] , \regIn[10][14] , 
        \regIn[10][13] , \regIn[10][12] , \regIn[10][11] , \regIn[10][10] , 
        \regIn[10][9] , \regIn[10][8] , \regIn[10][7] , \regIn[10][6] , 
        \regIn[10][5] , \regIn[10][4] , \regIn[10][3] , \regIn[10][2] , 
        \regIn[10][1] , \regIn[10][0] }), .clk(clk), .reset(n1273), .write(
        n1274), .dataOut({\regOut[10][15] , \regOut[10][14] , \regOut[10][13] , 
        \regOut[10][12] , \regOut[10][11] , \regOut[10][10] , \regOut[10][9] , 
        \regOut[10][8] , \regOut[10][7] , \regOut[10][6] , \regOut[10][5] , 
        \regOut[10][4] , \regOut[10][3] , \regOut[10][2] , \regOut[10][1] , 
        \regOut[10][0] }) );
  SingleReg_20 RegX_11 ( .data({\regIn[11][15] , \regIn[11][14] , 
        \regIn[11][13] , \regIn[11][12] , \regIn[11][11] , \regIn[11][10] , 
        \regIn[11][9] , \regIn[11][8] , \regIn[11][7] , \regIn[11][6] , 
        \regIn[11][5] , \regIn[11][4] , \regIn[11][3] , \regIn[11][2] , 
        \regIn[11][1] , \regIn[11][0] }), .clk(clk), .reset(n1273), .write(
        n1274), .dataOut({\regOut[11][15] , \regOut[11][14] , \regOut[11][13] , 
        \regOut[11][12] , \regOut[11][11] , \regOut[11][10] , \regOut[11][9] , 
        \regOut[11][8] , \regOut[11][7] , \regOut[11][6] , \regOut[11][5] , 
        \regOut[11][4] , \regOut[11][3] , \regOut[11][2] , \regOut[11][1] , 
        \regOut[11][0] }) );
  SingleReg_19 RegX_12 ( .data({\regIn[12][15] , \regIn[12][14] , 
        \regIn[12][13] , \regIn[12][12] , \regIn[12][11] , \regIn[12][10] , 
        \regIn[12][9] , \regIn[12][8] , \regIn[12][7] , \regIn[12][6] , 
        \regIn[12][5] , \regIn[12][4] , \regIn[12][3] , \regIn[12][2] , 
        \regIn[12][1] , \regIn[12][0] }), .clk(clk), .reset(n1273), .write(
        n1274), .dataOut({\regOut[12][15] , \regOut[12][14] , \regOut[12][13] , 
        \regOut[12][12] , \regOut[12][11] , \regOut[12][10] , \regOut[12][9] , 
        \regOut[12][8] , \regOut[12][7] , \regOut[12][6] , \regOut[12][5] , 
        \regOut[12][4] , \regOut[12][3] , \regOut[12][2] , \regOut[12][1] , 
        \regOut[12][0] }) );
  SingleReg_18 RegX_13 ( .data({\regIn[13][15] , \regIn[13][14] , 
        \regIn[13][13] , \regIn[13][12] , \regIn[13][11] , \regIn[13][10] , 
        \regIn[13][9] , \regIn[13][8] , \regIn[13][7] , \regIn[13][6] , 
        \regIn[13][5] , \regIn[13][4] , \regIn[13][3] , \regIn[13][2] , 
        \regIn[13][1] , \regIn[13][0] }), .clk(clk), .reset(n1273), .write(
        n1275), .dataOut({\regOut[13][15] , \regOut[13][14] , \regOut[13][13] , 
        \regOut[13][12] , \regOut[13][11] , \regOut[13][10] , \regOut[13][9] , 
        \regOut[13][8] , \regOut[13][7] , \regOut[13][6] , \regOut[13][5] , 
        \regOut[13][4] , \regOut[13][3] , \regOut[13][2] , \regOut[13][1] , 
        \regOut[13][0] }) );
  SingleReg_17 RegX_14 ( .data({\regIn[14][15] , \regIn[14][14] , 
        \regIn[14][13] , \regIn[14][12] , \regIn[14][11] , \regIn[14][10] , 
        \regIn[14][9] , \regIn[14][8] , \regIn[14][7] , \regIn[14][6] , 
        \regIn[14][5] , \regIn[14][4] , \regIn[14][3] , \regIn[14][2] , 
        \regIn[14][1] , \regIn[14][0] }), .clk(clk), .reset(n1273), .write(
        n1275), .dataOut({\regOut[14][15] , \regOut[14][14] , \regOut[14][13] , 
        \regOut[14][12] , \regOut[14][11] , \regOut[14][10] , \regOut[14][9] , 
        \regOut[14][8] , \regOut[14][7] , \regOut[14][6] , \regOut[14][5] , 
        \regOut[14][4] , \regOut[14][3] , \regOut[14][2] , \regOut[14][1] , 
        \regOut[14][0] }) );
  SingleReg_16 RegX_15 ( .data({\regIn[15][15] , \regIn[15][14] , 
        \regIn[15][13] , \regIn[15][12] , \regIn[15][11] , \regIn[15][10] , 
        \regIn[15][9] , \regIn[15][8] , \regIn[15][7] , \regIn[15][6] , 
        \regIn[15][5] , \regIn[15][4] , \regIn[15][3] , \regIn[15][2] , 
        \regIn[15][1] , \regIn[15][0] }), .clk(clk), .reset(n1273), .write(
        n1275), .dataOut({\regOut[15][15] , \regOut[15][14] , \regOut[15][13] , 
        \regOut[15][12] , \regOut[15][11] , \regOut[15][10] , \regOut[15][9] , 
        \regOut[15][8] , \regOut[15][7] , \regOut[15][6] , \regOut[15][5] , 
        \regOut[15][4] , \regOut[15][3] , \regOut[15][2] , \regOut[15][1] , 
        \regOut[15][0] }) );
  SingleReg_15 RegX_16 ( .data({\regIn[16][15] , \regIn[16][14] , 
        \regIn[16][13] , \regIn[16][12] , \regIn[16][11] , \regIn[16][10] , 
        \regIn[16][9] , \regIn[16][8] , \regIn[16][7] , \regIn[16][6] , 
        \regIn[16][5] , \regIn[16][4] , \regIn[16][3] , \regIn[16][2] , 
        \regIn[16][1] , \regIn[16][0] }), .clk(clk), .reset(n1273), .write(
        n1275), .dataOut({\regOut[16][15] , \regOut[16][14] , \regOut[16][13] , 
        \regOut[16][12] , \regOut[16][11] , \regOut[16][10] , \regOut[16][9] , 
        \regOut[16][8] , \regOut[16][7] , \regOut[16][6] , \regOut[16][5] , 
        \regOut[16][4] , \regOut[16][3] , \regOut[16][2] , \regOut[16][1] , 
        \regOut[16][0] }) );
  SingleReg_14 RegX_17 ( .data({\regIn[17][15] , \regIn[17][14] , 
        \regIn[17][13] , \regIn[17][12] , \regIn[17][11] , \regIn[17][10] , 
        \regIn[17][9] , \regIn[17][8] , \regIn[17][7] , \regIn[17][6] , 
        \regIn[17][5] , \regIn[17][4] , \regIn[17][3] , \regIn[17][2] , 
        \regIn[17][1] , \regIn[17][0] }), .clk(clk), .reset(n1273), .write(
        n1275), .dataOut({\regOut[17][15] , \regOut[17][14] , \regOut[17][13] , 
        \regOut[17][12] , \regOut[17][11] , \regOut[17][10] , \regOut[17][9] , 
        \regOut[17][8] , \regOut[17][7] , \regOut[17][6] , \regOut[17][5] , 
        \regOut[17][4] , \regOut[17][3] , \regOut[17][2] , \regOut[17][1] , 
        \regOut[17][0] }) );
  SingleReg_13 RegX_18 ( .data({\regIn[18][15] , \regIn[18][14] , 
        \regIn[18][13] , \regIn[18][12] , \regIn[18][11] , \regIn[18][10] , 
        \regIn[18][9] , \regIn[18][8] , \regIn[18][7] , \regIn[18][6] , 
        \regIn[18][5] , \regIn[18][4] , \regIn[18][3] , \regIn[18][2] , 
        \regIn[18][1] , \regIn[18][0] }), .clk(clk), .reset(n1273), .write(
        n1275), .dataOut({\regOut[18][15] , \regOut[18][14] , \regOut[18][13] , 
        \regOut[18][12] , \regOut[18][11] , \regOut[18][10] , \regOut[18][9] , 
        \regOut[18][8] , \regOut[18][7] , \regOut[18][6] , \regOut[18][5] , 
        \regOut[18][4] , \regOut[18][3] , \regOut[18][2] , \regOut[18][1] , 
        \regOut[18][0] }) );
  SingleReg_12 RegX_19 ( .data({\regIn[19][15] , \regIn[19][14] , 
        \regIn[19][13] , \regIn[19][12] , \regIn[19][11] , \regIn[19][10] , 
        \regIn[19][9] , \regIn[19][8] , \regIn[19][7] , \regIn[19][6] , 
        \regIn[19][5] , \regIn[19][4] , \regIn[19][3] , \regIn[19][2] , 
        \regIn[19][1] , \regIn[19][0] }), .clk(clk), .reset(n1273), .write(
        n1275), .dataOut({\regOut[19][15] , \regOut[19][14] , \regOut[19][13] , 
        \regOut[19][12] , \regOut[19][11] , \regOut[19][10] , \regOut[19][9] , 
        \regOut[19][8] , \regOut[19][7] , \regOut[19][6] , \regOut[19][5] , 
        \regOut[19][4] , \regOut[19][3] , \regOut[19][2] , \regOut[19][1] , 
        \regOut[19][0] }) );
  SingleReg_11 RegX_20 ( .data({\regIn[20][15] , \regIn[20][14] , 
        \regIn[20][13] , \regIn[20][12] , \regIn[20][11] , \regIn[20][10] , 
        \regIn[20][9] , \regIn[20][8] , \regIn[20][7] , \regIn[20][6] , 
        \regIn[20][5] , \regIn[20][4] , \regIn[20][3] , \regIn[20][2] , 
        \regIn[20][1] , \regIn[20][0] }), .clk(clk), .reset(n1273), .write(
        n1275), .dataOut({\regOut[20][15] , \regOut[20][14] , \regOut[20][13] , 
        \regOut[20][12] , \regOut[20][11] , \regOut[20][10] , \regOut[20][9] , 
        \regOut[20][8] , \regOut[20][7] , \regOut[20][6] , \regOut[20][5] , 
        \regOut[20][4] , \regOut[20][3] , \regOut[20][2] , \regOut[20][1] , 
        \regOut[20][0] }) );
  SingleReg_10 RegX_21 ( .data({\regIn[21][15] , \regIn[21][14] , 
        \regIn[21][13] , \regIn[21][12] , \regIn[21][11] , \regIn[21][10] , 
        \regIn[21][9] , \regIn[21][8] , \regIn[21][7] , \regIn[21][6] , 
        \regIn[21][5] , \regIn[21][4] , \regIn[21][3] , \regIn[21][2] , 
        \regIn[21][1] , \regIn[21][0] }), .clk(clk), .reset(n1273), .write(
        n1275), .dataOut({\regOut[21][15] , \regOut[21][14] , \regOut[21][13] , 
        \regOut[21][12] , \regOut[21][11] , \regOut[21][10] , \regOut[21][9] , 
        \regOut[21][8] , \regOut[21][7] , \regOut[21][6] , \regOut[21][5] , 
        \regOut[21][4] , \regOut[21][3] , \regOut[21][2] , \regOut[21][1] , 
        \regOut[21][0] }) );
  SingleReg_9 RegX_22 ( .data({\regIn[22][15] , \regIn[22][14] , 
        \regIn[22][13] , \regIn[22][12] , \regIn[22][11] , \regIn[22][10] , 
        \regIn[22][9] , \regIn[22][8] , \regIn[22][7] , \regIn[22][6] , 
        \regIn[22][5] , \regIn[22][4] , \regIn[22][3] , \regIn[22][2] , 
        \regIn[22][1] , \regIn[22][0] }), .clk(clk), .reset(n1273), .write(
        n1275), .dataOut({\regOut[22][15] , \regOut[22][14] , \regOut[22][13] , 
        \regOut[22][12] , \regOut[22][11] , \regOut[22][10] , \regOut[22][9] , 
        \regOut[22][8] , \regOut[22][7] , \regOut[22][6] , \regOut[22][5] , 
        \regOut[22][4] , \regOut[22][3] , \regOut[22][2] , \regOut[22][1] , 
        \regOut[22][0] }) );
  SingleReg_8 RegX_23 ( .data({\regIn[23][15] , \regIn[23][14] , 
        \regIn[23][13] , \regIn[23][12] , \regIn[23][11] , \regIn[23][10] , 
        \regIn[23][9] , \regIn[23][8] , \regIn[23][7] , \regIn[23][6] , 
        \regIn[23][5] , \regIn[23][4] , \regIn[23][3] , \regIn[23][2] , 
        \regIn[23][1] , \regIn[23][0] }), .clk(clk), .reset(n1273), .write(
        n1275), .dataOut({\regOut[23][15] , \regOut[23][14] , \regOut[23][13] , 
        \regOut[23][12] , \regOut[23][11] , \regOut[23][10] , \regOut[23][9] , 
        \regOut[23][8] , \regOut[23][7] , \regOut[23][6] , \regOut[23][5] , 
        \regOut[23][4] , \regOut[23][3] , \regOut[23][2] , \regOut[23][1] , 
        \regOut[23][0] }) );
  SingleReg_7 RegX_24 ( .data({\regIn[24][15] , \regIn[24][14] , 
        \regIn[24][13] , \regIn[24][12] , \regIn[24][11] , \regIn[24][10] , 
        \regIn[24][9] , \regIn[24][8] , \regIn[24][7] , \regIn[24][6] , 
        \regIn[24][5] , \regIn[24][4] , \regIn[24][3] , \regIn[24][2] , 
        \regIn[24][1] , \regIn[24][0] }), .clk(clk), .reset(n1273), .write(
        n1275), .dataOut({\regOut[24][15] , \regOut[24][14] , \regOut[24][13] , 
        \regOut[24][12] , \regOut[24][11] , \regOut[24][10] , \regOut[24][9] , 
        \regOut[24][8] , \regOut[24][7] , \regOut[24][6] , \regOut[24][5] , 
        \regOut[24][4] , \regOut[24][3] , \regOut[24][2] , \regOut[24][1] , 
        \regOut[24][0] }) );
  SingleReg_6 RegX_25 ( .data({\regIn[25][15] , \regIn[25][14] , 
        \regIn[25][13] , \regIn[25][12] , \regIn[25][11] , \regIn[25][10] , 
        \regIn[25][9] , \regIn[25][8] , \regIn[25][7] , \regIn[25][6] , 
        \regIn[25][5] , \regIn[25][4] , \regIn[25][3] , \regIn[25][2] , 
        \regIn[25][1] , \regIn[25][0] }), .clk(clk), .reset(n1273), .write(
        n1274), .dataOut({\regOut[25][15] , \regOut[25][14] , \regOut[25][13] , 
        \regOut[25][12] , \regOut[25][11] , \regOut[25][10] , \regOut[25][9] , 
        \regOut[25][8] , \regOut[25][7] , \regOut[25][6] , \regOut[25][5] , 
        \regOut[25][4] , \regOut[25][3] , \regOut[25][2] , \regOut[25][1] , 
        \regOut[25][0] }) );
  SingleReg_5 RegX_26 ( .data({\regIn[26][15] , \regIn[26][14] , 
        \regIn[26][13] , \regIn[26][12] , \regIn[26][11] , \regIn[26][10] , 
        \regIn[26][9] , \regIn[26][8] , \regIn[26][7] , \regIn[26][6] , 
        \regIn[26][5] , \regIn[26][4] , \regIn[26][3] , \regIn[26][2] , 
        \regIn[26][1] , \regIn[26][0] }), .clk(clk), .reset(n1273), .write(
        n1275), .dataOut({\regOut[26][15] , \regOut[26][14] , \regOut[26][13] , 
        \regOut[26][12] , \regOut[26][11] , \regOut[26][10] , \regOut[26][9] , 
        \regOut[26][8] , \regOut[26][7] , \regOut[26][6] , \regOut[26][5] , 
        \regOut[26][4] , \regOut[26][3] , \regOut[26][2] , \regOut[26][1] , 
        \regOut[26][0] }) );
  SingleReg_4 RegX_27 ( .data({\regIn[27][15] , \regIn[27][14] , 
        \regIn[27][13] , \regIn[27][12] , \regIn[27][11] , \regIn[27][10] , 
        \regIn[27][9] , \regIn[27][8] , \regIn[27][7] , \regIn[27][6] , 
        \regIn[27][5] , \regIn[27][4] , \regIn[27][3] , \regIn[27][2] , 
        \regIn[27][1] , \regIn[27][0] }), .clk(clk), .reset(n1273), .write(
        n1274), .dataOut({\regOut[27][15] , \regOut[27][14] , \regOut[27][13] , 
        \regOut[27][12] , \regOut[27][11] , \regOut[27][10] , \regOut[27][9] , 
        \regOut[27][8] , \regOut[27][7] , \regOut[27][6] , \regOut[27][5] , 
        \regOut[27][4] , \regOut[27][3] , \regOut[27][2] , \regOut[27][1] , 
        \regOut[27][0] }) );
  SingleReg_3 RegX_28 ( .data({\regIn[28][15] , \regIn[28][14] , 
        \regIn[28][13] , \regIn[28][12] , \regIn[28][11] , \regIn[28][10] , 
        \regIn[28][9] , \regIn[28][8] , \regIn[28][7] , \regIn[28][6] , 
        \regIn[28][5] , \regIn[28][4] , \regIn[28][3] , \regIn[28][2] , 
        \regIn[28][1] , \regIn[28][0] }), .clk(clk), .reset(n1273), .write(
        n1274), .dataOut({\regOut[28][15] , \regOut[28][14] , \regOut[28][13] , 
        \regOut[28][12] , \regOut[28][11] , \regOut[28][10] , \regOut[28][9] , 
        \regOut[28][8] , \regOut[28][7] , \regOut[28][6] , \regOut[28][5] , 
        \regOut[28][4] , \regOut[28][3] , \regOut[28][2] , \regOut[28][1] , 
        \regOut[28][0] }) );
  SingleReg_2 RegX_29 ( .data({\regIn[29][15] , \regIn[29][14] , 
        \regIn[29][13] , \regIn[29][12] , \regIn[29][11] , \regIn[29][10] , 
        \regIn[29][9] , \regIn[29][8] , \regIn[29][7] , \regIn[29][6] , 
        \regIn[29][5] , \regIn[29][4] , \regIn[29][3] , \regIn[29][2] , 
        \regIn[29][1] , \regIn[29][0] }), .clk(clk), .reset(n1273), .write(
        n1275), .dataOut({\regOut[29][15] , \regOut[29][14] , \regOut[29][13] , 
        \regOut[29][12] , \regOut[29][11] , \regOut[29][10] , \regOut[29][9] , 
        \regOut[29][8] , \regOut[29][7] , \regOut[29][6] , \regOut[29][5] , 
        \regOut[29][4] , \regOut[29][3] , \regOut[29][2] , \regOut[29][1] , 
        \regOut[29][0] }) );
  SingleReg_1 RegX_30 ( .data({\regIn[30][15] , \regIn[30][14] , 
        \regIn[30][13] , \regIn[30][12] , \regIn[30][11] , \regIn[30][10] , 
        \regIn[30][9] , \regIn[30][8] , \regIn[30][7] , \regIn[30][6] , 
        \regIn[30][5] , \regIn[30][4] , \regIn[30][3] , \regIn[30][2] , 
        \regIn[30][1] , \regIn[30][0] }), .clk(clk), .reset(n1273), .write(
        n1275), .dataOut({\regOut[30][15] , \regOut[30][14] , \regOut[30][13] , 
        \regOut[30][12] , \regOut[30][11] , \regOut[30][10] , \regOut[30][9] , 
        \regOut[30][8] , \regOut[30][7] , \regOut[30][6] , \regOut[30][5] , 
        \regOut[30][4] , \regOut[30][3] , \regOut[30][2] , \regOut[30][1] , 
        \regOut[30][0] }) );
  SingleReg_0 RegX_31 ( .data({\regIn[31][15] , \regIn[31][14] , 
        \regIn[31][13] , \regIn[31][12] , \regIn[31][11] , \regIn[31][10] , 
        \regIn[31][9] , \regIn[31][8] , \regIn[31][7] , \regIn[31][6] , 
        \regIn[31][5] , \regIn[31][4] , \regIn[31][3] , \regIn[31][2] , 
        \regIn[31][1] , \regIn[31][0] }), .clk(clk), .reset(n1273), .write(
        n1274), .dataOut({\regOut[31][15] , \regOut[31][14] , \regOut[31][13] , 
        \regOut[31][12] , \regOut[31][11] , \regOut[31][10] , \regOut[31][9] , 
        \regOut[31][8] , \regOut[31][7] , \regOut[31][6] , \regOut[31][5] , 
        \regOut[31][4] , \regOut[31][3] , \regOut[31][2] , \regOut[31][1] , 
        \regOut[31][0] }) );
  CLKBUF_X2 U1786 ( .A(write), .Z(n1274) );
  CLKBUF_X2 U1787 ( .A(write), .Z(n1275) );
  CLKBUF_X1 U1788 ( .A(addressA[1]), .Z(n1242) );
  CLKBUF_X1 U1789 ( .A(addressB[3]), .Z(n1243) );
  CLKBUF_X1 U1790 ( .A(addressA[2]), .Z(n1244) );
  CLKBUF_X1 U1791 ( .A(addressB[2]), .Z(n1245) );
  CLKBUF_X1 U1792 ( .A(addressA[3]), .Z(n1246) );
  CLKBUF_X1 U1793 ( .A(addressB[1]), .Z(n1247) );
  CLKBUF_X1 U1794 ( .A(addressA[4]), .Z(n1248) );
  CLKBUF_X1 U1795 ( .A(addressB[4]), .Z(n1249) );
  CLKBUF_X1 U1796 ( .A(addressA[0]), .Z(n1250) );
  CLKBUF_X1 U1797 ( .A(addressB[0]), .Z(n1251) );
  CLKBUF_X1 U1798 ( .A(dataIn[5]), .Z(n1252) );
  CLKBUF_X1 U1799 ( .A(dataIn[4]), .Z(n1253) );
  CLKBUF_X1 U1800 ( .A(dataIn[6]), .Z(n1254) );
  CLKBUF_X1 U1801 ( .A(dataIn[3]), .Z(n1255) );
  CLKBUF_X1 U1802 ( .A(dataIn[7]), .Z(n1256) );
  CLKBUF_X1 U1803 ( .A(dataIn[2]), .Z(n1257) );
  CLKBUF_X1 U1804 ( .A(dataIn[8]), .Z(n1258) );
  CLKBUF_X1 U1805 ( .A(dataIn[1]), .Z(n1259) );
  CLKBUF_X1 U1806 ( .A(dataIn[9]), .Z(n1260) );
  CLKBUF_X1 U1807 ( .A(dataIn[0]), .Z(n1261) );
  CLKBUF_X1 U1808 ( .A(dataIn[10]), .Z(n1262) );
  CLKBUF_X1 U1809 ( .A(addressIn[3]), .Z(n1263) );
  OR2_X1 U1810 ( .A1(n1263), .A2(N307), .ZN(N326) );
  OR2_X1 U1811 ( .A1(n1263), .A2(N307), .ZN(N302) );
  OR2_X1 U1812 ( .A1(n1263), .A2(N307), .ZN(N320) );
  OR2_X1 U1813 ( .A1(n1263), .A2(N307), .ZN(N296) );
  OR2_X1 U1814 ( .A1(n1263), .A2(N307), .ZN(N338) );
  OR2_X1 U1815 ( .A1(n1263), .A2(N307), .ZN(N314) );
  OR2_X1 U1816 ( .A1(n1263), .A2(N307), .ZN(N332) );
  INV_X1 U1817 ( .A(n1263), .ZN(N245) );
  OR2_X1 U1818 ( .A1(n1263), .A2(N307), .ZN(N308) );
  CLKBUF_X1 U1819 ( .A(dataIn[11]), .Z(n1264) );
  CLKBUF_X1 U1820 ( .A(addressIn[2]), .Z(n1265) );
  OR2_X1 U1821 ( .A1(n1265), .A2(N253), .ZN(N254) );
  OR2_X1 U1822 ( .A1(n1265), .A2(N350), .ZN(N351) );
  OR2_X1 U1823 ( .A1(n1265), .A2(N302), .ZN(N303) );
  OR2_X1 U1824 ( .A1(n1265), .A2(N202), .ZN(N203) );
  OR2_X1 U1825 ( .A1(n1265), .A2(N195), .ZN(N196) );
  OR2_X1 U1826 ( .A1(n1265), .A2(N247), .ZN(N248) );
  OR2_X1 U1827 ( .A1(n1265), .A2(N296), .ZN(N297) );
  OR2_X1 U1828 ( .A1(n1265), .A2(N344), .ZN(N345) );
  OR2_X1 U1829 ( .A1(n1265), .A2(N362), .ZN(N363) );
  OR2_X1 U1830 ( .A1(n1265), .A2(N215), .ZN(N216) );
  OR2_X1 U1831 ( .A1(n1265), .A2(N314), .ZN(N315) );
  OR2_X1 U1832 ( .A1(n1265), .A2(N265), .ZN(N266) );
  OR2_X1 U1833 ( .A1(n1265), .A2(N356), .ZN(N357) );
  OR2_X1 U1834 ( .A1(n1265), .A2(N209), .ZN(N210) );
  OR2_X1 U1835 ( .A1(n1265), .A2(N259), .ZN(N260) );
  OR2_X1 U1836 ( .A1(n1265), .A2(N308), .ZN(N309) );
  INV_X1 U1837 ( .A(n1265), .ZN(N220) );
  CLKBUF_X1 U1838 ( .A(dataIn[12]), .Z(n1266) );
  CLKBUF_X1 U1839 ( .A(addressIn[1]), .Z(n1267) );
  OR2_X1 U1840 ( .A1(n1267), .A2(N254), .ZN(N255) );
  OR2_X1 U1841 ( .A1(n1267), .A2(N351), .ZN(N352) );
  OR2_X1 U1842 ( .A1(n1267), .A2(N229), .ZN(N230) );
  OR2_X1 U1843 ( .A1(n1267), .A2(N303), .ZN(N304) );
  OR2_X1 U1844 ( .A1(n1267), .A2(N327), .ZN(N328) );
  OR2_X1 U1845 ( .A1(n1267), .A2(N203), .ZN(N204) );
  OR2_X1 U1846 ( .A1(n1267), .A2(N278), .ZN(N279) );
  OR2_X1 U1847 ( .A1(n1267), .A2(N196), .ZN(N197) );
  OR2_X1 U1848 ( .A1(n1267), .A2(N223), .ZN(N224) );
  OR2_X1 U1849 ( .A1(n1267), .A2(N272), .ZN(N273) );
  OR2_X1 U1850 ( .A1(n1267), .A2(N297), .ZN(N298) );
  OR2_X1 U1851 ( .A1(n1267), .A2(N321), .ZN(N322) );
  OR2_X1 U1852 ( .A1(n1267), .A2(N248), .ZN(N249) );
  OR2_X1 U1853 ( .A1(n1267), .A2(N345), .ZN(N346) );
  OR2_X1 U1854 ( .A1(n1267), .A2(N375), .ZN(N376) );
  OR2_X1 U1855 ( .A1(n1267), .A2(N369), .ZN(N370) );
  INV_X1 U1856 ( .A(n1267), .ZN(N207) );
  CLKBUF_X1 U1857 ( .A(dataIn[13]), .Z(n1268) );
  CLKBUF_X1 U1858 ( .A(addressIn[0]), .Z(n1269) );
  OR2_X1 U1859 ( .A1(n1269), .A2(N197), .ZN(N198) );
  OR2_X1 U1860 ( .A1(n1269), .A2(N382), .ZN(N383) );
  OR2_X1 U1861 ( .A1(n1269), .A2(N249), .ZN(N250) );
  OR2_X1 U1862 ( .A1(n1269), .A2(N346), .ZN(N347) );
  OR2_X1 U1863 ( .A1(n1269), .A2(N273), .ZN(N274) );
  OR2_X1 U1864 ( .A1(n1269), .A2(N224), .ZN(N225) );
  OR2_X1 U1865 ( .A1(n1269), .A2(N298), .ZN(N299) );
  OR2_X1 U1866 ( .A1(n1269), .A2(N322), .ZN(N323) );
  OR2_X1 U1867 ( .A1(n1269), .A2(N358), .ZN(N359) );
  OR2_X1 U1868 ( .A1(n1269), .A2(N370), .ZN(N371) );
  OR2_X1 U1869 ( .A1(n1269), .A2(N334), .ZN(N335) );
  OR2_X1 U1870 ( .A1(n1269), .A2(N211), .ZN(N212) );
  OR2_X1 U1871 ( .A1(n1269), .A2(N310), .ZN(N311) );
  OR2_X1 U1872 ( .A1(n1269), .A2(N261), .ZN(N262) );
  OR2_X1 U1873 ( .A1(n1269), .A2(N236), .ZN(N237) );
  OR2_X1 U1874 ( .A1(n1269), .A2(N285), .ZN(N286) );
  INV_X1 U1875 ( .A(n1269), .ZN(N200) );
  CLKBUF_X1 U1876 ( .A(dataIn[14]), .Z(n1270) );
  CLKBUF_X1 U1877 ( .A(N208), .Z(n1271) );
  OR2_X1 U1878 ( .A1(N245), .A2(n1271), .ZN(N253) );
  OR2_X1 U1879 ( .A1(N245), .A2(n1271), .ZN(N277) );
  OR2_X1 U1880 ( .A1(n1263), .A2(n1271), .ZN(N228) );
  OR2_X1 U1881 ( .A1(N245), .A2(n1271), .ZN(N271) );
  OR2_X1 U1882 ( .A1(n1263), .A2(n1271), .ZN(N202) );
  OR2_X1 U1883 ( .A1(n1263), .A2(n1271), .ZN(N222) );
  OR2_X1 U1884 ( .A1(N245), .A2(n1271), .ZN(N247) );
  OR2_X1 U1885 ( .A1(n1263), .A2(n1271), .ZN(N195) );
  OR2_X1 U1886 ( .A1(N245), .A2(n1271), .ZN(N289) );
  OR2_X1 U1887 ( .A1(n1263), .A2(n1271), .ZN(N240) );
  OR2_X1 U1888 ( .A1(N245), .A2(n1271), .ZN(N265) );
  OR2_X1 U1889 ( .A1(N245), .A2(n1271), .ZN(N283) );
  OR2_X1 U1890 ( .A1(n1263), .A2(n1271), .ZN(N215) );
  OR2_X1 U1891 ( .A1(n1263), .A2(n1271), .ZN(N234) );
  OR2_X1 U1892 ( .A1(N245), .A2(n1271), .ZN(N259) );
  OR2_X1 U1893 ( .A1(n1263), .A2(n1271), .ZN(N209) );
  INV_X1 U1894 ( .A(n1271), .ZN(N307) );
  CLKBUF_X1 U1895 ( .A(dataIn[15]), .Z(n1272) );
  CLKBUF_X2 U1896 ( .A(reset), .Z(n1273) );
endmodule

