module SingleReg_31 (
	data, 
	clk, 
	reset, 
	write, 
	dataOut, 
	FE_OFN1_write, 
	FE_OFN2_write, 
	FE_OFN18_write, 
	FE_OFN20_write, 
	FE_OFN22_write, 
	FE_OFN24_write, 
	FE_OFN29_write, 
	FE_OFN31_write, 
	clk__L2_N3, 
	clk__L2_N4, 
	clk__L2_N7, 
	clk__L2_N8, 
	VDD, 
	VSS);
   input [15:0] data;
   input clk;
   input reset;
   input write;
   output [15:0] dataOut;
   input FE_OFN1_write;
   input FE_OFN2_write;
   input FE_OFN18_write;
   input FE_OFN20_write;
   input FE_OFN22_write;
   input FE_OFN24_write;
   input FE_OFN29_write;
   input FE_OFN31_write;
   input clk__L2_N3;
   input clk__L2_N4;
   input clk__L2_N7;
   input clk__L2_N8;
   inout VDD;
   inout VSS;

   // Internal wires
   wire n1;
   wire n2;
   wire n3;
   wire n4;
   wire n5;
   wire n6;
   wire n7;
   wire n8;
   wire n9;
   wire n10;
   wire n11;
   wire n12;
   wire n13;
   wire n14;
   wire n15;
   wire n16;
   wire n17;
   wire n18;
   wire n19;
   wire n20;
   wire n21;
   wire n22;
   wire n23;
   wire n24;
   wire n25;
   wire n26;
   wire n27;
   wire n28;
   wire n29;
   wire n30;
   wire n31;
   wire n32;
   wire n33;
   wire n34;
   wire n35;
   wire n36;
   wire n37;
   wire n38;
   wire n39;
   wire n40;
   wire n41;
   wire n42;
   wire n43;
   wire n44;
   wire n45;
   wire n46;
   wire n47;
   wire n48;
   wire n49;

   // Module instantiations
   DFFR_X1 \Reg_reg[15]  (
	.RN(n48),
	.QN(n32),
	.Q(dataOut[15]),
	.D(n49),
	.CK(clk__L2_N7), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[14]  (
	.RN(n48),
	.QN(n31),
	.Q(dataOut[14]),
	.D(n47),
	.CK(clk__L2_N7), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[13]  (
	.RN(n48),
	.QN(n30),
	.Q(dataOut[13]),
	.D(n46),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[12]  (
	.RN(n48),
	.QN(n29),
	.Q(dataOut[12]),
	.D(n45),
	.CK(clk__L2_N7), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[11]  (
	.RN(n48),
	.QN(n28),
	.Q(dataOut[11]),
	.D(n44),
	.CK(clk__L2_N7), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[10]  (
	.RN(n48),
	.QN(n27),
	.Q(dataOut[10]),
	.D(n43),
	.CK(clk__L2_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[9]  (
	.RN(n48),
	.QN(n26),
	.Q(dataOut[9]),
	.D(n42),
	.CK(clk__L2_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[8]  (
	.RN(n48),
	.QN(n25),
	.Q(dataOut[8]),
	.D(n41),
	.CK(clk__L2_N7), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[7]  (
	.RN(n48),
	.QN(n24),
	.Q(dataOut[7]),
	.D(n40),
	.CK(clk__L2_N7), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[6]  (
	.RN(n48),
	.QN(n23),
	.Q(dataOut[6]),
	.D(n39),
	.CK(clk__L2_N7), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[5]  (
	.RN(n48),
	.QN(n22),
	.Q(dataOut[5]),
	.D(n38),
	.CK(clk__L2_N7), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[4]  (
	.RN(n48),
	.QN(n21),
	.Q(dataOut[4]),
	.D(n37),
	.CK(clk__L2_N8), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[3]  (
	.RN(n48),
	.QN(n20),
	.Q(dataOut[3]),
	.D(n36),
	.CK(clk__L2_N8), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[2]  (
	.RN(n48),
	.QN(n19),
	.Q(dataOut[2]),
	.D(n35),
	.CK(clk__L2_N7), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[1]  (
	.RN(n48),
	.QN(n18),
	.Q(dataOut[1]),
	.D(n34),
	.CK(clk__L2_N4), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[0]  (
	.RN(n48),
	.QN(n17),
	.Q(dataOut[0]),
	.D(n33),
	.CK(clk__L2_N8), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U2 (
	.ZN(n33),
	.B2(n17),
	.B1(FE_OFN18_write),
	.A(n1), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U3 (
	.ZN(n1),
	.A2(data[0]),
	.A1(FE_OFN18_write), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U4 (
	.ZN(n34),
	.B2(n18),
	.B1(FE_OFN1_write),
	.A(n2), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U5 (
	.ZN(n2),
	.A2(FE_OFN1_write),
	.A1(data[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U6 (
	.ZN(n35),
	.B2(n19),
	.B1(FE_OFN24_write),
	.A(n3), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U7 (
	.ZN(n3),
	.A2(FE_OFN24_write),
	.A1(data[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U8 (
	.ZN(n36),
	.B2(n20),
	.B1(FE_OFN1_write),
	.A(n4), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U9 (
	.ZN(n4),
	.A2(FE_OFN1_write),
	.A1(data[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U10 (
	.ZN(n37),
	.B2(n21),
	.B1(FE_OFN18_write),
	.A(n5), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U11 (
	.ZN(n5),
	.A2(FE_OFN18_write),
	.A1(data[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U12 (
	.ZN(n38),
	.B2(n22),
	.B1(FE_OFN22_write),
	.A(n6), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U13 (
	.ZN(n6),
	.A2(FE_OFN22_write),
	.A1(data[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U14 (
	.ZN(n39),
	.B2(n23),
	.B1(FE_OFN20_write),
	.A(n7), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U15 (
	.ZN(n7),
	.A2(FE_OFN20_write),
	.A1(data[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U16 (
	.ZN(n40),
	.B2(n24),
	.B1(write),
	.A(n8), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U17 (
	.ZN(n8),
	.A2(write),
	.A1(data[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U18 (
	.ZN(n41),
	.B2(n25),
	.B1(FE_OFN31_write),
	.A(n9), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U19 (
	.ZN(n9),
	.A2(FE_OFN31_write),
	.A1(data[8]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U20 (
	.ZN(n42),
	.B2(n26),
	.B1(FE_OFN29_write),
	.A(n10), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U21 (
	.ZN(n10),
	.A2(FE_OFN29_write),
	.A1(data[9]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U22 (
	.ZN(n43),
	.B2(n27),
	.B1(FE_OFN31_write),
	.A(n11), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U23 (
	.ZN(n11),
	.A2(FE_OFN31_write),
	.A1(data[10]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U24 (
	.ZN(n44),
	.B2(n28),
	.B1(FE_OFN20_write),
	.A(n12), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U25 (
	.ZN(n12),
	.A2(FE_OFN20_write),
	.A1(data[11]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U26 (
	.ZN(n45),
	.B2(n29),
	.B1(FE_OFN31_write),
	.A(n13), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U27 (
	.ZN(n13),
	.A2(FE_OFN31_write),
	.A1(data[12]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U28 (
	.ZN(n46),
	.B2(n30),
	.B1(FE_OFN2_write),
	.A(n14), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U29 (
	.ZN(n14),
	.A2(FE_OFN2_write),
	.A1(data[13]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U30 (
	.ZN(n47),
	.B2(n31),
	.B1(FE_OFN2_write),
	.A(n15), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U31 (
	.ZN(n15),
	.A2(FE_OFN2_write),
	.A1(data[14]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U32 (
	.ZN(n48),
	.A(reset), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U33 (
	.ZN(n49),
	.B2(n32),
	.B1(FE_OFN2_write),
	.A(n16), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U34 (
	.ZN(n16),
	.A2(FE_OFN2_write),
	.A1(data[15]), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module SingleReg_30 (
	data, 
	clk, 
	reset, 
	write, 
	dataOut, 
	FE_OFN1_write, 
	FE_OFN2_write, 
	FE_OFN18_write, 
	FE_OFN20_write, 
	FE_OFN22_write, 
	FE_OFN29_write, 
	FE_OFN31_write, 
	clk__L2_N3, 
	clk__L2_N4, 
	clk__L2_N7, 
	clk__L2_N8, 
	VDD, 
	VSS);
   input [15:0] data;
   input clk;
   input reset;
   input write;
   output [15:0] dataOut;
   input FE_OFN1_write;
   input FE_OFN2_write;
   input FE_OFN18_write;
   input FE_OFN20_write;
   input FE_OFN22_write;
   input FE_OFN29_write;
   input FE_OFN31_write;
   input clk__L2_N3;
   input clk__L2_N4;
   input clk__L2_N7;
   input clk__L2_N8;
   inout VDD;
   inout VSS;

   // Internal wires
   wire n53;
   wire n54;
   wire n55;
   wire n56;
   wire n57;
   wire n58;
   wire n59;
   wire n60;
   wire n61;
   wire n62;
   wire n63;
   wire n64;
   wire n65;
   wire n66;
   wire n67;
   wire n68;
   wire n69;
   wire n70;
   wire n71;
   wire n72;
   wire n73;
   wire n74;
   wire n75;
   wire n76;
   wire n77;
   wire n78;
   wire n79;
   wire n80;
   wire n81;
   wire n82;
   wire n83;
   wire n84;
   wire n85;
   wire n86;
   wire n87;
   wire n88;
   wire n89;
   wire n90;
   wire n91;
   wire n92;
   wire n93;
   wire n94;
   wire n95;
   wire n96;
   wire n97;
   wire n98;
   wire n99;
   wire n100;
   wire n101;

   // Module instantiations
   DFFR_X1 \Reg_reg[15]  (
	.RN(n54),
	.QN(n70),
	.Q(dataOut[15]),
	.D(n53),
	.CK(clk__L2_N7), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[14]  (
	.RN(n54),
	.QN(n71),
	.Q(dataOut[14]),
	.D(n55),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[13]  (
	.RN(n54),
	.QN(n72),
	.Q(dataOut[13]),
	.D(n56),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[12]  (
	.RN(n54),
	.QN(n73),
	.Q(dataOut[12]),
	.D(n57),
	.CK(clk__L2_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[11]  (
	.RN(n54),
	.QN(n74),
	.Q(dataOut[11]),
	.D(n58),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[10]  (
	.RN(n54),
	.QN(n75),
	.Q(dataOut[10]),
	.D(n59),
	.CK(clk__L2_N7), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[9]  (
	.RN(n54),
	.QN(n76),
	.Q(dataOut[9]),
	.D(n60),
	.CK(clk__L2_N7), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[8]  (
	.RN(n54),
	.QN(n77),
	.Q(dataOut[8]),
	.D(n61),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[7]  (
	.RN(n54),
	.QN(n78),
	.Q(dataOut[7]),
	.D(n62),
	.CK(clk__L2_N7), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[6]  (
	.RN(n54),
	.QN(n79),
	.Q(dataOut[6]),
	.D(n63),
	.CK(clk__L2_N7), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[5]  (
	.RN(n54),
	.QN(n80),
	.Q(dataOut[5]),
	.D(n64),
	.CK(clk__L2_N7), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[4]  (
	.RN(n54),
	.QN(n81),
	.Q(dataOut[4]),
	.D(n65),
	.CK(clk__L2_N8), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[3]  (
	.RN(n54),
	.QN(n82),
	.Q(dataOut[3]),
	.D(n66),
	.CK(clk__L2_N8), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[2]  (
	.RN(n54),
	.QN(n83),
	.Q(dataOut[2]),
	.D(n67),
	.CK(clk__L2_N4), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[1]  (
	.RN(n54),
	.QN(n84),
	.Q(dataOut[1]),
	.D(n68),
	.CK(clk__L2_N4), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[0]  (
	.RN(n54),
	.QN(n85),
	.Q(dataOut[0]),
	.D(n69),
	.CK(clk__L2_N8), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U2 (
	.ZN(n69),
	.B2(n85),
	.B1(FE_OFN18_write),
	.A(n101), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U3 (
	.ZN(n101),
	.A2(data[0]),
	.A1(FE_OFN18_write), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U4 (
	.ZN(n68),
	.B2(n84),
	.B1(FE_OFN18_write),
	.A(n100), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U5 (
	.ZN(n100),
	.A2(FE_OFN18_write),
	.A1(data[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U6 (
	.ZN(n67),
	.B2(n83),
	.B1(FE_OFN18_write),
	.A(n99), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U7 (
	.ZN(n99),
	.A2(FE_OFN18_write),
	.A1(data[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U8 (
	.ZN(n66),
	.B2(n82),
	.B1(FE_OFN18_write),
	.A(n98), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U9 (
	.ZN(n98),
	.A2(FE_OFN18_write),
	.A1(data[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U10 (
	.ZN(n65),
	.B2(n81),
	.B1(write),
	.A(n97), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U11 (
	.ZN(n97),
	.A2(FE_OFN1_write),
	.A1(data[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U12 (
	.ZN(n64),
	.B2(n80),
	.B1(FE_OFN1_write),
	.A(n96), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U13 (
	.ZN(n96),
	.A2(FE_OFN22_write),
	.A1(data[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U14 (
	.ZN(n63),
	.B2(n79),
	.B1(FE_OFN20_write),
	.A(n95), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U15 (
	.ZN(n95),
	.A2(FE_OFN20_write),
	.A1(data[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U16 (
	.ZN(n62),
	.B2(n78),
	.B1(FE_OFN29_write),
	.A(n94), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U17 (
	.ZN(n94),
	.A2(FE_OFN29_write),
	.A1(data[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U18 (
	.ZN(n61),
	.B2(n77),
	.B1(FE_OFN2_write),
	.A(n93), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U19 (
	.ZN(n93),
	.A2(FE_OFN2_write),
	.A1(data[8]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U20 (
	.ZN(n60),
	.B2(n76),
	.B1(FE_OFN22_write),
	.A(n92), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U21 (
	.ZN(n92),
	.A2(FE_OFN22_write),
	.A1(data[9]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U22 (
	.ZN(n59),
	.B2(n75),
	.B1(FE_OFN29_write),
	.A(n91), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U23 (
	.ZN(n91),
	.A2(FE_OFN31_write),
	.A1(data[10]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U24 (
	.ZN(n58),
	.B2(n74),
	.B1(FE_OFN31_write),
	.A(n90), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U25 (
	.ZN(n90),
	.A2(FE_OFN31_write),
	.A1(data[11]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U26 (
	.ZN(n57),
	.B2(n73),
	.B1(FE_OFN31_write),
	.A(n89), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U27 (
	.ZN(n89),
	.A2(FE_OFN31_write),
	.A1(data[12]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U28 (
	.ZN(n56),
	.B2(n72),
	.B1(FE_OFN2_write),
	.A(n88), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U29 (
	.ZN(n88),
	.A2(FE_OFN2_write),
	.A1(data[13]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U30 (
	.ZN(n55),
	.B2(n71),
	.B1(FE_OFN2_write),
	.A(n87), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U31 (
	.ZN(n87),
	.A2(FE_OFN2_write),
	.A1(data[14]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X2 U32 (
	.ZN(n54),
	.A(reset), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U33 (
	.ZN(n53),
	.B2(n70),
	.B1(FE_OFN20_write),
	.A(n86), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U34 (
	.ZN(n86),
	.A2(FE_OFN20_write),
	.A1(data[15]), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module SingleReg_29 (
	data, 
	clk, 
	reset, 
	write, 
	dataOut, 
	FE_OFN0_write, 
	FE_OFN15_write, 
	FE_OFN16_write, 
	FE_OFN17_write, 
	clk__L2_N8, 
	VDD, 
	VSS);
   input [15:0] data;
   input clk;
   input reset;
   input write;
   output [15:0] dataOut;
   input FE_OFN0_write;
   input FE_OFN15_write;
   input FE_OFN16_write;
   input FE_OFN17_write;
   input clk__L2_N8;
   inout VDD;
   inout VSS;

   // Internal wires
   wire n53;
   wire n54;
   wire n55;
   wire n56;
   wire n57;
   wire n58;
   wire n59;
   wire n60;
   wire n61;
   wire n62;
   wire n63;
   wire n64;
   wire n65;
   wire n66;
   wire n67;
   wire n68;
   wire n69;
   wire n70;
   wire n71;
   wire n72;
   wire n73;
   wire n74;
   wire n75;
   wire n76;
   wire n77;
   wire n78;
   wire n79;
   wire n80;
   wire n81;
   wire n82;
   wire n83;
   wire n84;
   wire n85;
   wire n86;
   wire n87;
   wire n88;
   wire n89;
   wire n90;
   wire n91;
   wire n92;
   wire n93;
   wire n94;
   wire n95;
   wire n96;
   wire n97;
   wire n98;
   wire n99;
   wire n100;
   wire n101;

   // Module instantiations
   DFFR_X1 \Reg_reg[15]  (
	.RN(n54),
	.QN(n70),
	.Q(dataOut[15]),
	.D(n53),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[14]  (
	.RN(n54),
	.QN(n71),
	.Q(dataOut[14]),
	.D(n55),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[13]  (
	.RN(n54),
	.QN(n72),
	.Q(dataOut[13]),
	.D(n56),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[12]  (
	.RN(n54),
	.QN(n73),
	.Q(dataOut[12]),
	.D(n57),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[11]  (
	.RN(n54),
	.QN(n74),
	.Q(dataOut[11]),
	.D(n58),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[10]  (
	.RN(n54),
	.QN(n75),
	.Q(dataOut[10]),
	.D(n59),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[9]  (
	.RN(n54),
	.QN(n76),
	.Q(dataOut[9]),
	.D(n60),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[8]  (
	.RN(n54),
	.QN(n77),
	.Q(dataOut[8]),
	.D(n61),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[7]  (
	.RN(n54),
	.QN(n78),
	.Q(dataOut[7]),
	.D(n62),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[6]  (
	.RN(n54),
	.QN(n79),
	.Q(dataOut[6]),
	.D(n63),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[5]  (
	.RN(n54),
	.QN(n80),
	.Q(dataOut[5]),
	.D(n64),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[4]  (
	.RN(n54),
	.QN(n81),
	.Q(dataOut[4]),
	.D(n65),
	.CK(clk__L2_N8), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[3]  (
	.RN(n54),
	.QN(n82),
	.Q(dataOut[3]),
	.D(n66),
	.CK(clk__L2_N8), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[2]  (
	.RN(n54),
	.QN(n83),
	.Q(dataOut[2]),
	.D(n67),
	.CK(clk__L2_N8), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[1]  (
	.RN(n54),
	.QN(n84),
	.Q(dataOut[1]),
	.D(n68),
	.CK(clk__L2_N8), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[0]  (
	.RN(n54),
	.QN(n85),
	.Q(dataOut[0]),
	.D(n69),
	.CK(clk__L2_N8), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U2 (
	.ZN(n69),
	.B2(n85),
	.B1(FE_OFN17_write),
	.A(n101), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U3 (
	.ZN(n101),
	.A2(data[0]),
	.A1(FE_OFN17_write), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U4 (
	.ZN(n68),
	.B2(n84),
	.B1(FE_OFN17_write),
	.A(n100), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U5 (
	.ZN(n100),
	.A2(FE_OFN17_write),
	.A1(data[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U6 (
	.ZN(n67),
	.B2(n83),
	.B1(FE_OFN17_write),
	.A(n99), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U7 (
	.ZN(n99),
	.A2(FE_OFN17_write),
	.A1(data[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U8 (
	.ZN(n66),
	.B2(n82),
	.B1(write),
	.A(n98), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U9 (
	.ZN(n98),
	.A2(write),
	.A1(data[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U10 (
	.ZN(n65),
	.B2(n81),
	.B1(FE_OFN16_write),
	.A(n97), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U11 (
	.ZN(n97),
	.A2(FE_OFN0_write),
	.A1(data[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U12 (
	.ZN(n64),
	.B2(n80),
	.B1(write),
	.A(n96), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U13 (
	.ZN(n96),
	.A2(write),
	.A1(data[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U14 (
	.ZN(n63),
	.B2(n79),
	.B1(FE_OFN16_write),
	.A(n95), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U15 (
	.ZN(n95),
	.A2(FE_OFN16_write),
	.A1(data[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U16 (
	.ZN(n62),
	.B2(n78),
	.B1(FE_OFN16_write),
	.A(n94), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U17 (
	.ZN(n94),
	.A2(FE_OFN15_write),
	.A1(data[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U18 (
	.ZN(n61),
	.B2(n77),
	.B1(FE_OFN16_write),
	.A(n93), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U19 (
	.ZN(n93),
	.A2(FE_OFN16_write),
	.A1(data[8]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U20 (
	.ZN(n60),
	.B2(n76),
	.B1(FE_OFN16_write),
	.A(n92), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U21 (
	.ZN(n92),
	.A2(FE_OFN16_write),
	.A1(data[9]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U22 (
	.ZN(n59),
	.B2(n75),
	.B1(FE_OFN16_write),
	.A(n91), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U23 (
	.ZN(n91),
	.A2(FE_OFN16_write),
	.A1(data[10]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U24 (
	.ZN(n58),
	.B2(n74),
	.B1(FE_OFN16_write),
	.A(n90), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U25 (
	.ZN(n90),
	.A2(FE_OFN16_write),
	.A1(data[11]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U26 (
	.ZN(n57),
	.B2(n73),
	.B1(FE_OFN16_write),
	.A(n89), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U27 (
	.ZN(n89),
	.A2(FE_OFN16_write),
	.A1(data[12]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U28 (
	.ZN(n56),
	.B2(n72),
	.B1(FE_OFN16_write),
	.A(n88), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U29 (
	.ZN(n88),
	.A2(FE_OFN16_write),
	.A1(data[13]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U30 (
	.ZN(n55),
	.B2(n71),
	.B1(FE_OFN16_write),
	.A(n87), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U31 (
	.ZN(n87),
	.A2(FE_OFN16_write),
	.A1(data[14]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U32 (
	.ZN(n54),
	.A(reset), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U33 (
	.ZN(n53),
	.B2(n70),
	.B1(FE_OFN16_write),
	.A(n86), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U34 (
	.ZN(n86),
	.A2(FE_OFN16_write),
	.A1(data[15]), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module SingleReg_28 (
	data, 
	clk, 
	reset, 
	write, 
	dataOut, 
	FE_OFN0_write, 
	FE_OFN17_write, 
	FE_OFN18_write, 
	FE_OFN20_write, 
	clk__L2_N8, 
	VDD, 
	VSS);
   input [15:0] data;
   input clk;
   input reset;
   input write;
   output [15:0] dataOut;
   input FE_OFN0_write;
   input FE_OFN17_write;
   input FE_OFN18_write;
   input FE_OFN20_write;
   input clk__L2_N8;
   inout VDD;
   inout VSS;

   // Internal wires
   wire FE_OFN19_write;
   wire n53;
   wire n54;
   wire n55;
   wire n56;
   wire n57;
   wire n58;
   wire n59;
   wire n60;
   wire n61;
   wire n62;
   wire n63;
   wire n64;
   wire n65;
   wire n66;
   wire n67;
   wire n68;
   wire n69;
   wire n70;
   wire n71;
   wire n72;
   wire n73;
   wire n74;
   wire n75;
   wire n76;
   wire n77;
   wire n78;
   wire n79;
   wire n80;
   wire n81;
   wire n82;
   wire n83;
   wire n84;
   wire n85;
   wire n86;
   wire n87;
   wire n88;
   wire n89;
   wire n90;
   wire n91;
   wire n92;
   wire n93;
   wire n94;
   wire n95;
   wire n96;
   wire n97;
   wire n98;
   wire n99;
   wire n100;
   wire n101;

   // Module instantiations
   CLKBUF_X1 FE_OFC19_write (
	.Z(FE_OFN19_write),
	.A(FE_OFN18_write), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[15]  (
	.RN(n54),
	.QN(n70),
	.Q(dataOut[15]),
	.D(n53),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[14]  (
	.RN(n54),
	.QN(n71),
	.Q(dataOut[14]),
	.D(n55),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[13]  (
	.RN(n54),
	.QN(n72),
	.Q(dataOut[13]),
	.D(n56),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[12]  (
	.RN(n54),
	.QN(n73),
	.Q(dataOut[12]),
	.D(n57),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[11]  (
	.RN(n54),
	.QN(n74),
	.Q(dataOut[11]),
	.D(n58),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[10]  (
	.RN(n54),
	.QN(n75),
	.Q(dataOut[10]),
	.D(n59),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[9]  (
	.RN(n54),
	.QN(n76),
	.Q(dataOut[9]),
	.D(n60),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[8]  (
	.RN(n54),
	.QN(n77),
	.Q(dataOut[8]),
	.D(n61),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[7]  (
	.RN(n54),
	.QN(n78),
	.Q(dataOut[7]),
	.D(n62),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[6]  (
	.RN(n54),
	.QN(n79),
	.Q(dataOut[6]),
	.D(n63),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[5]  (
	.RN(n54),
	.QN(n80),
	.Q(dataOut[5]),
	.D(n64),
	.CK(clk__L2_N8), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[4]  (
	.RN(n54),
	.QN(n81),
	.Q(dataOut[4]),
	.D(n65),
	.CK(clk__L2_N8), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[3]  (
	.RN(n54),
	.QN(n82),
	.Q(dataOut[3]),
	.D(n66),
	.CK(clk__L2_N8), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[2]  (
	.RN(n54),
	.QN(n83),
	.Q(dataOut[2]),
	.D(n67),
	.CK(clk__L2_N8), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[1]  (
	.RN(n54),
	.QN(n84),
	.Q(dataOut[1]),
	.D(n68),
	.CK(clk__L2_N8), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[0]  (
	.RN(n54),
	.QN(n85),
	.Q(dataOut[0]),
	.D(n69),
	.CK(clk__L2_N8), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U2 (
	.ZN(n69),
	.B2(n85),
	.B1(FE_OFN19_write),
	.A(n101), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U3 (
	.ZN(n101),
	.A2(data[0]),
	.A1(FE_OFN19_write), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U4 (
	.ZN(n68),
	.B2(n84),
	.B1(FE_OFN19_write),
	.A(n100), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U5 (
	.ZN(n100),
	.A2(FE_OFN19_write),
	.A1(data[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U6 (
	.ZN(n67),
	.B2(n83),
	.B1(FE_OFN18_write),
	.A(n99), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U7 (
	.ZN(n99),
	.A2(FE_OFN18_write),
	.A1(data[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U8 (
	.ZN(n66),
	.B2(n82),
	.B1(FE_OFN17_write),
	.A(n98), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U9 (
	.ZN(n98),
	.A2(FE_OFN19_write),
	.A1(data[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U10 (
	.ZN(n65),
	.B2(n81),
	.B1(FE_OFN0_write),
	.A(n97), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U11 (
	.ZN(n97),
	.A2(FE_OFN0_write),
	.A1(data[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U12 (
	.ZN(n64),
	.B2(n80),
	.B1(FE_OFN0_write),
	.A(n96), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U13 (
	.ZN(n96),
	.A2(FE_OFN0_write),
	.A1(data[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U14 (
	.ZN(n63),
	.B2(n79),
	.B1(write),
	.A(n95), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U15 (
	.ZN(n95),
	.A2(FE_OFN0_write),
	.A1(data[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U16 (
	.ZN(n62),
	.B2(n78),
	.B1(FE_OFN0_write),
	.A(n94), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U17 (
	.ZN(n94),
	.A2(FE_OFN0_write),
	.A1(data[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U18 (
	.ZN(n61),
	.B2(n77),
	.B1(write),
	.A(n93), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U19 (
	.ZN(n93),
	.A2(write),
	.A1(data[8]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U20 (
	.ZN(n60),
	.B2(n76),
	.B1(FE_OFN0_write),
	.A(n92), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U21 (
	.ZN(n92),
	.A2(FE_OFN20_write),
	.A1(data[9]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U22 (
	.ZN(n59),
	.B2(n75),
	.B1(write),
	.A(n91), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U23 (
	.ZN(n91),
	.A2(write),
	.A1(data[10]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U24 (
	.ZN(n58),
	.B2(n74),
	.B1(FE_OFN20_write),
	.A(n90), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U25 (
	.ZN(n90),
	.A2(FE_OFN20_write),
	.A1(data[11]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U26 (
	.ZN(n57),
	.B2(n73),
	.B1(write),
	.A(n89), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U27 (
	.ZN(n89),
	.A2(write),
	.A1(data[12]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U28 (
	.ZN(n56),
	.B2(n72),
	.B1(FE_OFN20_write),
	.A(n88), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U29 (
	.ZN(n88),
	.A2(FE_OFN20_write),
	.A1(data[13]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U30 (
	.ZN(n55),
	.B2(n71),
	.B1(write),
	.A(n87), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U31 (
	.ZN(n87),
	.A2(write),
	.A1(data[14]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U32 (
	.ZN(n54),
	.A(reset), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U33 (
	.ZN(n53),
	.B2(n70),
	.B1(write),
	.A(n86), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U34 (
	.ZN(n86),
	.A2(write),
	.A1(data[15]), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module SingleReg_27 (
	data, 
	clk, 
	reset, 
	write, 
	dataOut, 
	FE_OFN5_write, 
	FE_OFN6_write, 
	FE_OFN32_write, 
	FE_OFN36_write, 
	FE_OFN44_write, 
	clk__L2_N2, 
	clk__L2_N3, 
	VDD, 
	VSS);
   input [15:0] data;
   input clk;
   input reset;
   input write;
   output [15:0] dataOut;
   input FE_OFN5_write;
   input FE_OFN6_write;
   input FE_OFN32_write;
   input FE_OFN36_write;
   input FE_OFN44_write;
   input clk__L2_N2;
   input clk__L2_N3;
   inout VDD;
   inout VSS;

   // Internal wires
   wire n53;
   wire n54;
   wire n55;
   wire n56;
   wire n57;
   wire n58;
   wire n59;
   wire n60;
   wire n61;
   wire n62;
   wire n63;
   wire n64;
   wire n65;
   wire n66;
   wire n67;
   wire n68;
   wire n69;
   wire n70;
   wire n71;
   wire n72;
   wire n73;
   wire n74;
   wire n75;
   wire n76;
   wire n77;
   wire n78;
   wire n79;
   wire n80;
   wire n81;
   wire n82;
   wire n83;
   wire n84;
   wire n85;
   wire n86;
   wire n87;
   wire n88;
   wire n89;
   wire n90;
   wire n91;
   wire n92;
   wire n93;
   wire n94;
   wire n95;
   wire n96;
   wire n97;
   wire n98;
   wire n99;
   wire n100;
   wire n101;

   // Module instantiations
   DFFR_X1 \Reg_reg[15]  (
	.RN(n54),
	.QN(n70),
	.Q(dataOut[15]),
	.D(n53),
	.CK(clk__L2_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[14]  (
	.RN(n54),
	.QN(n71),
	.Q(dataOut[14]),
	.D(n55),
	.CK(clk__L2_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[13]  (
	.RN(n54),
	.QN(n72),
	.Q(dataOut[13]),
	.D(n56),
	.CK(clk__L2_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[12]  (
	.RN(n54),
	.QN(n73),
	.Q(dataOut[12]),
	.D(n57),
	.CK(clk__L2_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[11]  (
	.RN(n54),
	.QN(n74),
	.Q(dataOut[11]),
	.D(n58),
	.CK(clk__L2_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[10]  (
	.RN(n54),
	.QN(n75),
	.Q(dataOut[10]),
	.D(n59),
	.CK(clk__L2_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[9]  (
	.RN(n54),
	.QN(n76),
	.Q(dataOut[9]),
	.D(n60),
	.CK(clk__L2_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[8]  (
	.RN(n54),
	.QN(n77),
	.Q(dataOut[8]),
	.D(n61),
	.CK(clk__L2_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[7]  (
	.RN(n54),
	.QN(n78),
	.Q(dataOut[7]),
	.D(n62),
	.CK(clk__L2_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[6]  (
	.RN(n54),
	.QN(n79),
	.Q(dataOut[6]),
	.D(n63),
	.CK(clk__L2_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[5]  (
	.RN(n54),
	.QN(n80),
	.Q(dataOut[5]),
	.D(n64),
	.CK(clk__L2_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[4]  (
	.RN(n54),
	.QN(n81),
	.Q(dataOut[4]),
	.D(n65),
	.CK(clk__L2_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[3]  (
	.RN(n54),
	.QN(n82),
	.Q(dataOut[3]),
	.D(n66),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[2]  (
	.RN(n54),
	.QN(n83),
	.Q(dataOut[2]),
	.D(n67),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[1]  (
	.RN(n54),
	.QN(n84),
	.Q(dataOut[1]),
	.D(n68),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[0]  (
	.RN(n54),
	.QN(n85),
	.Q(dataOut[0]),
	.D(n69),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U2 (
	.ZN(n69),
	.B2(n85),
	.B1(FE_OFN5_write),
	.A(n101), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U3 (
	.ZN(n101),
	.A2(data[0]),
	.A1(FE_OFN5_write), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U4 (
	.ZN(n68),
	.B2(n84),
	.B1(FE_OFN5_write),
	.A(n100), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U5 (
	.ZN(n100),
	.A2(FE_OFN5_write),
	.A1(data[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U6 (
	.ZN(n67),
	.B2(n83),
	.B1(FE_OFN5_write),
	.A(n99), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U7 (
	.ZN(n99),
	.A2(FE_OFN5_write),
	.A1(data[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U8 (
	.ZN(n66),
	.B2(n82),
	.B1(FE_OFN5_write),
	.A(n98), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U9 (
	.ZN(n98),
	.A2(FE_OFN5_write),
	.A1(data[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U10 (
	.ZN(n65),
	.B2(n81),
	.B1(FE_OFN32_write),
	.A(n97), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U11 (
	.ZN(n97),
	.A2(FE_OFN32_write),
	.A1(data[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U12 (
	.ZN(n64),
	.B2(n80),
	.B1(write),
	.A(n96), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U13 (
	.ZN(n96),
	.A2(write),
	.A1(data[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U14 (
	.ZN(n63),
	.B2(n79),
	.B1(FE_OFN32_write),
	.A(n95), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U15 (
	.ZN(n95),
	.A2(FE_OFN32_write),
	.A1(data[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U16 (
	.ZN(n62),
	.B2(n78),
	.B1(write),
	.A(n94), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U17 (
	.ZN(n94),
	.A2(write),
	.A1(data[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U18 (
	.ZN(n61),
	.B2(n77),
	.B1(FE_OFN6_write),
	.A(n93), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U19 (
	.ZN(n93),
	.A2(FE_OFN6_write),
	.A1(data[8]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U20 (
	.ZN(n60),
	.B2(n76),
	.B1(write),
	.A(n92), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U21 (
	.ZN(n92),
	.A2(write),
	.A1(data[9]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U22 (
	.ZN(n59),
	.B2(n75),
	.B1(FE_OFN44_write),
	.A(n91), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U23 (
	.ZN(n91),
	.A2(FE_OFN44_write),
	.A1(data[10]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U24 (
	.ZN(n58),
	.B2(n74),
	.B1(FE_OFN32_write),
	.A(n90), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U25 (
	.ZN(n90),
	.A2(FE_OFN32_write),
	.A1(data[11]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U26 (
	.ZN(n57),
	.B2(n73),
	.B1(FE_OFN32_write),
	.A(n89), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U27 (
	.ZN(n89),
	.A2(FE_OFN32_write),
	.A1(data[12]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U28 (
	.ZN(n56),
	.B2(n72),
	.B1(FE_OFN44_write),
	.A(n88), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U29 (
	.ZN(n88),
	.A2(FE_OFN44_write),
	.A1(data[13]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U30 (
	.ZN(n55),
	.B2(n71),
	.B1(FE_OFN44_write),
	.A(n87), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U31 (
	.ZN(n87),
	.A2(FE_OFN44_write),
	.A1(data[14]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X2 U32 (
	.ZN(n54),
	.A(reset), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U33 (
	.ZN(n53),
	.B2(n70),
	.B1(FE_OFN44_write),
	.A(n86), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U34 (
	.ZN(n86),
	.A2(FE_OFN44_write),
	.A1(data[15]), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module SingleReg_26 (
	data, 
	clk, 
	reset, 
	write, 
	dataOut, 
	FE_OFN5_write, 
	FE_OFN6_write, 
	FE_OFN32_write, 
	FE_OFN36_write, 
	clk__L2_N2, 
	clk__L2_N3, 
	VDD, 
	VSS);
   input [15:0] data;
   input clk;
   input reset;
   input write;
   output [15:0] dataOut;
   input FE_OFN5_write;
   input FE_OFN6_write;
   input FE_OFN32_write;
   input FE_OFN36_write;
   input clk__L2_N2;
   input clk__L2_N3;
   inout VDD;
   inout VSS;

   // Internal wires
   wire n53;
   wire n54;
   wire n55;
   wire n56;
   wire n57;
   wire n58;
   wire n59;
   wire n60;
   wire n61;
   wire n62;
   wire n63;
   wire n64;
   wire n65;
   wire n66;
   wire n67;
   wire n68;
   wire n69;
   wire n70;
   wire n71;
   wire n72;
   wire n73;
   wire n74;
   wire n75;
   wire n76;
   wire n77;
   wire n78;
   wire n79;
   wire n80;
   wire n81;
   wire n82;
   wire n83;
   wire n84;
   wire n85;
   wire n86;
   wire n87;
   wire n88;
   wire n89;
   wire n90;
   wire n91;
   wire n92;
   wire n93;
   wire n94;
   wire n95;
   wire n96;
   wire n97;
   wire n98;
   wire n99;
   wire n100;
   wire n101;

   // Module instantiations
   DFFR_X1 \Reg_reg[15]  (
	.RN(n54),
	.QN(n70),
	.Q(dataOut[15]),
	.D(n53),
	.CK(clk__L2_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[14]  (
	.RN(n54),
	.QN(n71),
	.Q(dataOut[14]),
	.D(n55),
	.CK(clk__L2_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[13]  (
	.RN(n54),
	.QN(n72),
	.Q(dataOut[13]),
	.D(n56),
	.CK(clk__L2_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[12]  (
	.RN(n54),
	.QN(n73),
	.Q(dataOut[12]),
	.D(n57),
	.CK(clk__L2_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[11]  (
	.RN(n54),
	.QN(n74),
	.Q(dataOut[11]),
	.D(n58),
	.CK(clk__L2_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[10]  (
	.RN(n54),
	.QN(n75),
	.Q(dataOut[10]),
	.D(n59),
	.CK(clk__L2_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[9]  (
	.RN(n54),
	.QN(n76),
	.Q(dataOut[9]),
	.D(n60),
	.CK(clk__L2_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[8]  (
	.RN(n54),
	.QN(n77),
	.Q(dataOut[8]),
	.D(n61),
	.CK(clk__L2_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[7]  (
	.RN(n54),
	.QN(n78),
	.Q(dataOut[7]),
	.D(n62),
	.CK(clk__L2_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[6]  (
	.RN(n54),
	.QN(n79),
	.Q(dataOut[6]),
	.D(n63),
	.CK(clk__L2_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[5]  (
	.RN(n54),
	.QN(n80),
	.Q(dataOut[5]),
	.D(n64),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[4]  (
	.RN(n54),
	.QN(n81),
	.Q(dataOut[4]),
	.D(n65),
	.CK(clk__L2_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[3]  (
	.RN(n54),
	.QN(n82),
	.Q(dataOut[3]),
	.D(n66),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[2]  (
	.RN(n54),
	.QN(n83),
	.Q(dataOut[2]),
	.D(n67),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[1]  (
	.RN(n54),
	.QN(n84),
	.Q(dataOut[1]),
	.D(n68),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[0]  (
	.RN(n54),
	.QN(n85),
	.Q(dataOut[0]),
	.D(n69),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U2 (
	.ZN(n69),
	.B2(n85),
	.B1(FE_OFN5_write),
	.A(n101), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U3 (
	.ZN(n101),
	.A2(data[0]),
	.A1(FE_OFN5_write), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U4 (
	.ZN(n68),
	.B2(n84),
	.B1(FE_OFN5_write),
	.A(n100), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U5 (
	.ZN(n100),
	.A2(FE_OFN5_write),
	.A1(data[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U6 (
	.ZN(n67),
	.B2(n83),
	.B1(FE_OFN5_write),
	.A(n99), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U7 (
	.ZN(n99),
	.A2(FE_OFN5_write),
	.A1(data[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U8 (
	.ZN(n66),
	.B2(n82),
	.B1(FE_OFN5_write),
	.A(n98), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U9 (
	.ZN(n98),
	.A2(FE_OFN5_write),
	.A1(data[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U10 (
	.ZN(n65),
	.B2(n81),
	.B1(write),
	.A(n97), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U11 (
	.ZN(n97),
	.A2(write),
	.A1(data[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U12 (
	.ZN(n64),
	.B2(n80),
	.B1(write),
	.A(n96), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U13 (
	.ZN(n96),
	.A2(write),
	.A1(data[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U14 (
	.ZN(n63),
	.B2(n79),
	.B1(write),
	.A(n95), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U15 (
	.ZN(n95),
	.A2(write),
	.A1(data[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U16 (
	.ZN(n62),
	.B2(n78),
	.B1(write),
	.A(n94), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U17 (
	.ZN(n94),
	.A2(write),
	.A1(data[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U18 (
	.ZN(n61),
	.B2(n77),
	.B1(FE_OFN32_write),
	.A(n93), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U19 (
	.ZN(n93),
	.A2(FE_OFN32_write),
	.A1(data[8]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U20 (
	.ZN(n60),
	.B2(n76),
	.B1(FE_OFN32_write),
	.A(n92), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U21 (
	.ZN(n92),
	.A2(FE_OFN32_write),
	.A1(data[9]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U22 (
	.ZN(n59),
	.B2(n75),
	.B1(FE_OFN6_write),
	.A(n91), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U23 (
	.ZN(n91),
	.A2(FE_OFN6_write),
	.A1(data[10]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U24 (
	.ZN(n58),
	.B2(n74),
	.B1(FE_OFN32_write),
	.A(n90), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U25 (
	.ZN(n90),
	.A2(FE_OFN32_write),
	.A1(data[11]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U26 (
	.ZN(n57),
	.B2(n73),
	.B1(FE_OFN32_write),
	.A(n89), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U27 (
	.ZN(n89),
	.A2(FE_OFN32_write),
	.A1(data[12]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U28 (
	.ZN(n56),
	.B2(n72),
	.B1(FE_OFN6_write),
	.A(n88), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U29 (
	.ZN(n88),
	.A2(FE_OFN6_write),
	.A1(data[13]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U30 (
	.ZN(n55),
	.B2(n71),
	.B1(FE_OFN6_write),
	.A(n87), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U31 (
	.ZN(n87),
	.A2(FE_OFN6_write),
	.A1(data[14]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X2 U32 (
	.ZN(n54),
	.A(reset), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U33 (
	.ZN(n53),
	.B2(n70),
	.B1(FE_OFN32_write),
	.A(n86), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U34 (
	.ZN(n86),
	.A2(FE_OFN32_write),
	.A1(data[15]), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module SingleReg_25 (
	data, 
	clk, 
	reset, 
	write, 
	dataOut, 
	FE_OFN2_write, 
	FE_OFN6_write, 
	FE_OFN25_write, 
	FE_OFN31_write, 
	FE_OFN32_write, 
	FE_OFN41_write, 
	clk__L2_N2, 
	clk__L2_N3, 
	clk__L2_N4, 
	VDD, 
	VSS);
   input [15:0] data;
   input clk;
   input reset;
   input write;
   output [15:0] dataOut;
   input FE_OFN2_write;
   input FE_OFN6_write;
   input FE_OFN25_write;
   input FE_OFN31_write;
   input FE_OFN32_write;
   input FE_OFN41_write;
   input clk__L2_N2;
   input clk__L2_N3;
   input clk__L2_N4;
   inout VDD;
   inout VSS;

   // Internal wires
   wire n53;
   wire n54;
   wire n55;
   wire n56;
   wire n57;
   wire n58;
   wire n59;
   wire n60;
   wire n61;
   wire n62;
   wire n63;
   wire n64;
   wire n65;
   wire n66;
   wire n67;
   wire n68;
   wire n69;
   wire n70;
   wire n71;
   wire n72;
   wire n73;
   wire n74;
   wire n75;
   wire n76;
   wire n77;
   wire n78;
   wire n79;
   wire n80;
   wire n81;
   wire n82;
   wire n83;
   wire n84;
   wire n85;
   wire n86;
   wire n87;
   wire n88;
   wire n89;
   wire n90;
   wire n91;
   wire n92;
   wire n93;
   wire n94;
   wire n95;
   wire n96;
   wire n97;
   wire n98;
   wire n99;
   wire n100;
   wire n101;

   // Module instantiations
   DFFR_X1 \Reg_reg[15]  (
	.RN(n54),
	.QN(n70),
	.Q(dataOut[15]),
	.D(n53),
	.CK(clk__L2_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[14]  (
	.RN(n54),
	.QN(n71),
	.Q(dataOut[14]),
	.D(n55),
	.CK(clk__L2_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[13]  (
	.RN(n54),
	.QN(n72),
	.Q(dataOut[13]),
	.D(n56),
	.CK(clk__L2_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[12]  (
	.RN(n54),
	.QN(n73),
	.Q(dataOut[12]),
	.D(n57),
	.CK(clk__L2_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[11]  (
	.RN(n54),
	.QN(n74),
	.Q(dataOut[11]),
	.D(n58),
	.CK(clk__L2_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[10]  (
	.RN(n54),
	.QN(n75),
	.Q(dataOut[10]),
	.D(n59),
	.CK(clk__L2_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[9]  (
	.RN(n54),
	.QN(n76),
	.Q(dataOut[9]),
	.D(n60),
	.CK(clk__L2_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[8]  (
	.RN(n54),
	.QN(n77),
	.Q(dataOut[8]),
	.D(n61),
	.CK(clk__L2_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[7]  (
	.RN(n54),
	.QN(n78),
	.Q(dataOut[7]),
	.D(n62),
	.CK(clk__L2_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[6]  (
	.RN(n54),
	.QN(n79),
	.Q(dataOut[6]),
	.D(n63),
	.CK(clk__L2_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[5]  (
	.RN(n54),
	.QN(n80),
	.Q(dataOut[5]),
	.D(n64),
	.CK(clk__L2_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[4]  (
	.RN(n54),
	.QN(n81),
	.Q(dataOut[4]),
	.D(n65),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[3]  (
	.RN(n54),
	.QN(n82),
	.Q(dataOut[3]),
	.D(n66),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[2]  (
	.RN(n54),
	.QN(n83),
	.Q(dataOut[2]),
	.D(n67),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[1]  (
	.RN(n54),
	.QN(n84),
	.Q(dataOut[1]),
	.D(n68),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[0]  (
	.RN(n54),
	.QN(n85),
	.Q(dataOut[0]),
	.D(n69),
	.CK(clk__L2_N4), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U2 (
	.ZN(n69),
	.B2(n85),
	.B1(FE_OFN25_write),
	.A(n101), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U3 (
	.ZN(n101),
	.A2(data[0]),
	.A1(FE_OFN25_write), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U4 (
	.ZN(n68),
	.B2(n84),
	.B1(FE_OFN25_write),
	.A(n100), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U5 (
	.ZN(n100),
	.A2(FE_OFN25_write),
	.A1(data[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U6 (
	.ZN(n67),
	.B2(n83),
	.B1(FE_OFN25_write),
	.A(n99), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U7 (
	.ZN(n99),
	.A2(FE_OFN25_write),
	.A1(data[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U8 (
	.ZN(n66),
	.B2(n82),
	.B1(FE_OFN25_write),
	.A(n98), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U9 (
	.ZN(n98),
	.A2(FE_OFN25_write),
	.A1(data[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U10 (
	.ZN(n65),
	.B2(n81),
	.B1(write),
	.A(n97), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U11 (
	.ZN(n97),
	.A2(write),
	.A1(data[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U12 (
	.ZN(n64),
	.B2(n80),
	.B1(write),
	.A(n96), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U13 (
	.ZN(n96),
	.A2(write),
	.A1(data[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U14 (
	.ZN(n63),
	.B2(n79),
	.B1(FE_OFN31_write),
	.A(n95), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U15 (
	.ZN(n95),
	.A2(FE_OFN31_write),
	.A1(data[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U16 (
	.ZN(n62),
	.B2(n78),
	.B1(write),
	.A(n94), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U17 (
	.ZN(n94),
	.A2(write),
	.A1(data[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U18 (
	.ZN(n61),
	.B2(n77),
	.B1(FE_OFN6_write),
	.A(n93), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U19 (
	.ZN(n93),
	.A2(FE_OFN6_write),
	.A1(data[8]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U20 (
	.ZN(n60),
	.B2(n76),
	.B1(FE_OFN2_write),
	.A(n92), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U21 (
	.ZN(n92),
	.A2(FE_OFN2_write),
	.A1(data[9]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U22 (
	.ZN(n59),
	.B2(n75),
	.B1(FE_OFN31_write),
	.A(n91), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U23 (
	.ZN(n91),
	.A2(FE_OFN31_write),
	.A1(data[10]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U24 (
	.ZN(n58),
	.B2(n74),
	.B1(FE_OFN31_write),
	.A(n90), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U25 (
	.ZN(n90),
	.A2(FE_OFN31_write),
	.A1(data[11]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U26 (
	.ZN(n57),
	.B2(n73),
	.B1(FE_OFN41_write),
	.A(n89), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U27 (
	.ZN(n89),
	.A2(FE_OFN41_write),
	.A1(data[12]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U28 (
	.ZN(n56),
	.B2(n72),
	.B1(FE_OFN32_write),
	.A(n88), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U29 (
	.ZN(n88),
	.A2(FE_OFN32_write),
	.A1(data[13]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U30 (
	.ZN(n55),
	.B2(n71),
	.B1(FE_OFN41_write),
	.A(n87), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U31 (
	.ZN(n87),
	.A2(FE_OFN41_write),
	.A1(data[14]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U32 (
	.ZN(n54),
	.A(reset), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U33 (
	.ZN(n53),
	.B2(n70),
	.B1(FE_OFN41_write),
	.A(n86), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U34 (
	.ZN(n86),
	.A2(FE_OFN41_write),
	.A1(data[15]), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module SingleReg_24 (
	data, 
	clk, 
	reset, 
	write, 
	dataOut, 
	FE_OFN2_write, 
	FE_OFN24_write, 
	FE_OFN25_write, 
	FE_OFN31_write, 
	clk__L2_N2, 
	clk__L2_N3, 
	clk__L2_N4, 
	VDD, 
	VSS);
   input [15:0] data;
   input clk;
   input reset;
   input write;
   output [15:0] dataOut;
   input FE_OFN2_write;
   input FE_OFN24_write;
   input FE_OFN25_write;
   input FE_OFN31_write;
   input clk__L2_N2;
   input clk__L2_N3;
   input clk__L2_N4;
   inout VDD;
   inout VSS;

   // Internal wires
   wire n53;
   wire n54;
   wire n55;
   wire n56;
   wire n57;
   wire n58;
   wire n59;
   wire n60;
   wire n61;
   wire n62;
   wire n63;
   wire n64;
   wire n65;
   wire n66;
   wire n67;
   wire n68;
   wire n69;
   wire n70;
   wire n71;
   wire n72;
   wire n73;
   wire n74;
   wire n75;
   wire n76;
   wire n77;
   wire n78;
   wire n79;
   wire n80;
   wire n81;
   wire n82;
   wire n83;
   wire n84;
   wire n85;
   wire n86;
   wire n87;
   wire n88;
   wire n89;
   wire n90;
   wire n91;
   wire n92;
   wire n93;
   wire n94;
   wire n95;
   wire n96;
   wire n97;
   wire n98;
   wire n99;
   wire n100;
   wire n101;

   // Module instantiations
   DFFR_X1 \Reg_reg[15]  (
	.RN(n54),
	.QN(n70),
	.Q(dataOut[15]),
	.D(n53),
	.CK(clk__L2_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[14]  (
	.RN(n54),
	.QN(n71),
	.Q(dataOut[14]),
	.D(n55),
	.CK(clk__L2_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[13]  (
	.RN(n54),
	.QN(n72),
	.Q(dataOut[13]),
	.D(n56),
	.CK(clk__L2_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[12]  (
	.RN(n54),
	.QN(n73),
	.Q(dataOut[12]),
	.D(n57),
	.CK(clk__L2_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[11]  (
	.RN(n54),
	.QN(n74),
	.Q(dataOut[11]),
	.D(n58),
	.CK(clk__L2_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[10]  (
	.RN(n54),
	.QN(n75),
	.Q(dataOut[10]),
	.D(n59),
	.CK(clk__L2_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[9]  (
	.RN(n54),
	.QN(n76),
	.Q(dataOut[9]),
	.D(n60),
	.CK(clk__L2_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[8]  (
	.RN(n54),
	.QN(n77),
	.Q(dataOut[8]),
	.D(n61),
	.CK(clk__L2_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[7]  (
	.RN(n54),
	.QN(n78),
	.Q(dataOut[7]),
	.D(n62),
	.CK(clk__L2_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[6]  (
	.RN(n54),
	.QN(n79),
	.Q(dataOut[6]),
	.D(n63),
	.CK(clk__L2_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[5]  (
	.RN(n54),
	.QN(n80),
	.Q(dataOut[5]),
	.D(n64),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[4]  (
	.RN(n54),
	.QN(n81),
	.Q(dataOut[4]),
	.D(n65),
	.CK(clk__L2_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[3]  (
	.RN(n54),
	.QN(n82),
	.Q(dataOut[3]),
	.D(n66),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[2]  (
	.RN(n54),
	.QN(n83),
	.Q(dataOut[2]),
	.D(n67),
	.CK(clk__L2_N4), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[1]  (
	.RN(n54),
	.QN(n84),
	.Q(dataOut[1]),
	.D(n68),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[0]  (
	.RN(n54),
	.QN(n85),
	.Q(dataOut[0]),
	.D(n69),
	.CK(clk__L2_N4), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U2 (
	.ZN(n69),
	.B2(n85),
	.B1(FE_OFN24_write),
	.A(n101), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U3 (
	.ZN(n101),
	.A2(data[0]),
	.A1(FE_OFN24_write), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U4 (
	.ZN(n68),
	.B2(n84),
	.B1(FE_OFN25_write),
	.A(n100), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U5 (
	.ZN(n100),
	.A2(FE_OFN25_write),
	.A1(data[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U6 (
	.ZN(n67),
	.B2(n83),
	.B1(write),
	.A(n99), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U7 (
	.ZN(n99),
	.A2(write),
	.A1(data[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U8 (
	.ZN(n66),
	.B2(n82),
	.B1(write),
	.A(n98), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U9 (
	.ZN(n98),
	.A2(FE_OFN25_write),
	.A1(data[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U10 (
	.ZN(n65),
	.B2(n81),
	.B1(write),
	.A(n97), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U11 (
	.ZN(n97),
	.A2(write),
	.A1(data[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U12 (
	.ZN(n64),
	.B2(n80),
	.B1(write),
	.A(n96), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U13 (
	.ZN(n96),
	.A2(write),
	.A1(data[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U14 (
	.ZN(n63),
	.B2(n79),
	.B1(FE_OFN31_write),
	.A(n95), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U15 (
	.ZN(n95),
	.A2(FE_OFN31_write),
	.A1(data[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U16 (
	.ZN(n62),
	.B2(n78),
	.B1(write),
	.A(n94), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U17 (
	.ZN(n94),
	.A2(write),
	.A1(data[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U18 (
	.ZN(n61),
	.B2(n77),
	.B1(FE_OFN2_write),
	.A(n93), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U19 (
	.ZN(n93),
	.A2(FE_OFN2_write),
	.A1(data[8]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U20 (
	.ZN(n60),
	.B2(n76),
	.B1(write),
	.A(n92), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U21 (
	.ZN(n92),
	.A2(write),
	.A1(data[9]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U22 (
	.ZN(n59),
	.B2(n75),
	.B1(FE_OFN31_write),
	.A(n91), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U23 (
	.ZN(n91),
	.A2(FE_OFN31_write),
	.A1(data[10]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U24 (
	.ZN(n58),
	.B2(n74),
	.B1(FE_OFN31_write),
	.A(n90), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U25 (
	.ZN(n90),
	.A2(FE_OFN31_write),
	.A1(data[11]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U26 (
	.ZN(n57),
	.B2(n73),
	.B1(FE_OFN2_write),
	.A(n89), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U27 (
	.ZN(n89),
	.A2(FE_OFN2_write),
	.A1(data[12]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U28 (
	.ZN(n56),
	.B2(n72),
	.B1(FE_OFN2_write),
	.A(n88), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U29 (
	.ZN(n88),
	.A2(FE_OFN2_write),
	.A1(data[13]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U30 (
	.ZN(n55),
	.B2(n71),
	.B1(FE_OFN2_write),
	.A(n87), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U31 (
	.ZN(n87),
	.A2(FE_OFN2_write),
	.A1(data[14]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U32 (
	.ZN(n54),
	.A(reset), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U33 (
	.ZN(n53),
	.B2(n70),
	.B1(FE_OFN2_write),
	.A(n86), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U34 (
	.ZN(n86),
	.A2(FE_OFN2_write),
	.A1(data[15]), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module SingleReg_23 (
	data, 
	clk, 
	reset, 
	write, 
	dataOut, 
	FE_OFN4_write, 
	FE_OFN6_write, 
	FE_OFN34_write, 
	FE_OFN43_write, 
	clk__L2_N12, 
	clk__L2_N2, 
	clk__L2_N3, 
	VDD, 
	VSS);
   input [15:0] data;
   input clk;
   input reset;
   input write;
   output [15:0] dataOut;
   input FE_OFN4_write;
   input FE_OFN6_write;
   input FE_OFN34_write;
   input FE_OFN43_write;
   input clk__L2_N12;
   input clk__L2_N2;
   input clk__L2_N3;
   inout VDD;
   inout VSS;

   // Internal wires
   wire FE_OFN33_write;
   wire n53;
   wire n54;
   wire n55;
   wire n56;
   wire n57;
   wire n58;
   wire n59;
   wire n60;
   wire n61;
   wire n62;
   wire n63;
   wire n64;
   wire n65;
   wire n66;
   wire n67;
   wire n68;
   wire n69;
   wire n70;
   wire n71;
   wire n72;
   wire n73;
   wire n74;
   wire n75;
   wire n76;
   wire n77;
   wire n78;
   wire n79;
   wire n80;
   wire n81;
   wire n82;
   wire n83;
   wire n84;
   wire n85;
   wire n86;
   wire n87;
   wire n88;
   wire n89;
   wire n90;
   wire n91;
   wire n92;
   wire n93;
   wire n94;
   wire n95;
   wire n96;
   wire n97;
   wire n98;
   wire n99;
   wire n100;
   wire n101;

   // Module instantiations
   CLKBUF_X1 FE_OFC33_write (
	.Z(FE_OFN33_write),
	.A(FE_OFN4_write), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[15]  (
	.RN(n54),
	.QN(n70),
	.Q(dataOut[15]),
	.D(n53),
	.CK(clk__L2_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[14]  (
	.RN(n54),
	.QN(n71),
	.Q(dataOut[14]),
	.D(n55),
	.CK(clk__L2_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[13]  (
	.RN(n54),
	.QN(n72),
	.Q(dataOut[13]),
	.D(n56),
	.CK(clk__L2_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[12]  (
	.RN(n54),
	.QN(n73),
	.Q(dataOut[12]),
	.D(n57),
	.CK(clk__L2_N12), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[11]  (
	.RN(n54),
	.QN(n74),
	.Q(dataOut[11]),
	.D(n58),
	.CK(clk__L2_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[10]  (
	.RN(n54),
	.QN(n75),
	.Q(dataOut[10]),
	.D(n59),
	.CK(clk__L2_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[9]  (
	.RN(n54),
	.QN(n76),
	.Q(dataOut[9]),
	.D(n60),
	.CK(clk__L2_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[8]  (
	.RN(n54),
	.QN(n77),
	.Q(dataOut[8]),
	.D(n61),
	.CK(clk__L2_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[7]  (
	.RN(n54),
	.QN(n78),
	.Q(dataOut[7]),
	.D(n62),
	.CK(clk__L2_N12), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[6]  (
	.RN(n54),
	.QN(n79),
	.Q(dataOut[6]),
	.D(n63),
	.CK(clk__L2_N12), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[5]  (
	.RN(n54),
	.QN(n80),
	.Q(dataOut[5]),
	.D(n64),
	.CK(clk__L2_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[4]  (
	.RN(n54),
	.QN(n81),
	.Q(dataOut[4]),
	.D(n65),
	.CK(clk__L2_N12), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[3]  (
	.RN(n54),
	.QN(n82),
	.Q(dataOut[3]),
	.D(n66),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[2]  (
	.RN(n54),
	.QN(n83),
	.Q(dataOut[2]),
	.D(n67),
	.CK(clk__L2_N12), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[1]  (
	.RN(n54),
	.QN(n84),
	.Q(dataOut[1]),
	.D(n68),
	.CK(clk__L2_N12), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[0]  (
	.RN(n54),
	.QN(n85),
	.Q(dataOut[0]),
	.D(n69),
	.CK(clk__L2_N12), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U2 (
	.ZN(n69),
	.B2(n85),
	.B1(FE_OFN43_write),
	.A(n101), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U3 (
	.ZN(n101),
	.A2(data[0]),
	.A1(FE_OFN43_write), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U4 (
	.ZN(n68),
	.B2(n84),
	.B1(FE_OFN43_write),
	.A(n100), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U5 (
	.ZN(n100),
	.A2(FE_OFN43_write),
	.A1(data[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U6 (
	.ZN(n67),
	.B2(n83),
	.B1(FE_OFN33_write),
	.A(n99), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U7 (
	.ZN(n99),
	.A2(FE_OFN33_write),
	.A1(data[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U8 (
	.ZN(n66),
	.B2(n82),
	.B1(FE_OFN33_write),
	.A(n98), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U9 (
	.ZN(n98),
	.A2(FE_OFN33_write),
	.A1(data[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U10 (
	.ZN(n65),
	.B2(n81),
	.B1(FE_OFN4_write),
	.A(n97), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U11 (
	.ZN(n97),
	.A2(FE_OFN4_write),
	.A1(data[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U12 (
	.ZN(n64),
	.B2(n80),
	.B1(FE_OFN33_write),
	.A(n96), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U13 (
	.ZN(n96),
	.A2(FE_OFN33_write),
	.A1(data[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U14 (
	.ZN(n63),
	.B2(n79),
	.B1(FE_OFN34_write),
	.A(n95), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U15 (
	.ZN(n95),
	.A2(FE_OFN34_write),
	.A1(data[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U16 (
	.ZN(n62),
	.B2(n78),
	.B1(FE_OFN4_write),
	.A(n94), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U17 (
	.ZN(n94),
	.A2(FE_OFN4_write),
	.A1(data[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U18 (
	.ZN(n61),
	.B2(n77),
	.B1(FE_OFN6_write),
	.A(n93), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U19 (
	.ZN(n93),
	.A2(FE_OFN6_write),
	.A1(data[8]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U20 (
	.ZN(n60),
	.B2(n76),
	.B1(FE_OFN34_write),
	.A(n92), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U21 (
	.ZN(n92),
	.A2(FE_OFN34_write),
	.A1(data[9]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U22 (
	.ZN(n59),
	.B2(n75),
	.B1(write),
	.A(n91), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U23 (
	.ZN(n91),
	.A2(write),
	.A1(data[10]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U24 (
	.ZN(n58),
	.B2(n74),
	.B1(write),
	.A(n90), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U25 (
	.ZN(n90),
	.A2(write),
	.A1(data[11]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U26 (
	.ZN(n57),
	.B2(n73),
	.B1(FE_OFN34_write),
	.A(n89), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U27 (
	.ZN(n89),
	.A2(FE_OFN34_write),
	.A1(data[12]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U28 (
	.ZN(n56),
	.B2(n72),
	.B1(FE_OFN6_write),
	.A(n88), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U29 (
	.ZN(n88),
	.A2(FE_OFN6_write),
	.A1(data[13]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U30 (
	.ZN(n55),
	.B2(n71),
	.B1(FE_OFN6_write),
	.A(n87), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U31 (
	.ZN(n87),
	.A2(FE_OFN6_write),
	.A1(data[14]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U32 (
	.ZN(n54),
	.A(reset), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U33 (
	.ZN(n53),
	.B2(n70),
	.B1(FE_OFN6_write),
	.A(n86), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U34 (
	.ZN(n86),
	.A2(FE_OFN6_write),
	.A1(data[15]), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module SingleReg_22 (
	data, 
	clk, 
	reset, 
	write, 
	dataOut, 
	FE_OFN5_write, 
	FE_OFN6_write, 
	FE_OFN34_write, 
	FE_OFN47_write, 
	clk__L2_N12, 
	clk__L2_N2, 
	clk__L2_N3, 
	VDD, 
	VSS);
   input [15:0] data;
   input clk;
   input reset;
   input write;
   output [15:0] dataOut;
   input FE_OFN5_write;
   input FE_OFN6_write;
   input FE_OFN34_write;
   input FE_OFN47_write;
   input clk__L2_N12;
   input clk__L2_N2;
   input clk__L2_N3;
   inout VDD;
   inout VSS;

   // Internal wires
   wire n53;
   wire n54;
   wire n55;
   wire n56;
   wire n57;
   wire n58;
   wire n59;
   wire n60;
   wire n61;
   wire n62;
   wire n63;
   wire n64;
   wire n65;
   wire n66;
   wire n67;
   wire n68;
   wire n69;
   wire n70;
   wire n71;
   wire n72;
   wire n73;
   wire n74;
   wire n75;
   wire n76;
   wire n77;
   wire n78;
   wire n79;
   wire n80;
   wire n81;
   wire n82;
   wire n83;
   wire n84;
   wire n85;
   wire n86;
   wire n87;
   wire n88;
   wire n89;
   wire n90;
   wire n91;
   wire n92;
   wire n93;
   wire n94;
   wire n95;
   wire n96;
   wire n97;
   wire n98;
   wire n99;
   wire n100;
   wire n101;

   // Module instantiations
   DFFR_X1 \Reg_reg[15]  (
	.RN(n54),
	.QN(n70),
	.Q(dataOut[15]),
	.D(n53),
	.CK(clk__L2_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[14]  (
	.RN(n54),
	.QN(n71),
	.Q(dataOut[14]),
	.D(n55),
	.CK(clk__L2_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[13]  (
	.RN(n54),
	.QN(n72),
	.Q(dataOut[13]),
	.D(n56),
	.CK(clk__L2_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[12]  (
	.RN(n54),
	.QN(n73),
	.Q(dataOut[12]),
	.D(n57),
	.CK(clk__L2_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[11]  (
	.RN(n54),
	.QN(n74),
	.Q(dataOut[11]),
	.D(n58),
	.CK(clk__L2_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[10]  (
	.RN(n54),
	.QN(n75),
	.Q(dataOut[10]),
	.D(n59),
	.CK(clk__L2_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[9]  (
	.RN(n54),
	.QN(n76),
	.Q(dataOut[9]),
	.D(n60),
	.CK(clk__L2_N12), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[8]  (
	.RN(n54),
	.QN(n77),
	.Q(dataOut[8]),
	.D(n61),
	.CK(clk__L2_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[7]  (
	.RN(n54),
	.QN(n78),
	.Q(dataOut[7]),
	.D(n62),
	.CK(clk__L2_N12), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[6]  (
	.RN(n54),
	.QN(n79),
	.Q(dataOut[6]),
	.D(n63),
	.CK(clk__L2_N12), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[5]  (
	.RN(n54),
	.QN(n80),
	.Q(dataOut[5]),
	.D(n64),
	.CK(clk__L2_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[4]  (
	.RN(n54),
	.QN(n81),
	.Q(dataOut[4]),
	.D(n65),
	.CK(clk__L2_N12), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[3]  (
	.RN(n54),
	.QN(n82),
	.Q(dataOut[3]),
	.D(n66),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[2]  (
	.RN(n54),
	.QN(n83),
	.Q(dataOut[2]),
	.D(n67),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[1]  (
	.RN(n54),
	.QN(n84),
	.Q(dataOut[1]),
	.D(n68),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[0]  (
	.RN(n54),
	.QN(n85),
	.Q(dataOut[0]),
	.D(n69),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U2 (
	.ZN(n69),
	.B2(n85),
	.B1(FE_OFN47_write),
	.A(n101), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U3 (
	.ZN(n101),
	.A2(data[0]),
	.A1(FE_OFN5_write), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U4 (
	.ZN(n68),
	.B2(n84),
	.B1(FE_OFN47_write),
	.A(n100), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U5 (
	.ZN(n100),
	.A2(FE_OFN47_write),
	.A1(data[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U6 (
	.ZN(n67),
	.B2(n83),
	.B1(FE_OFN5_write),
	.A(n99), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U7 (
	.ZN(n99),
	.A2(FE_OFN5_write),
	.A1(data[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U8 (
	.ZN(n66),
	.B2(n82),
	.B1(FE_OFN5_write),
	.A(n98), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U9 (
	.ZN(n98),
	.A2(FE_OFN5_write),
	.A1(data[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U10 (
	.ZN(n65),
	.B2(n81),
	.B1(write),
	.A(n97), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U11 (
	.ZN(n97),
	.A2(write),
	.A1(data[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U12 (
	.ZN(n64),
	.B2(n80),
	.B1(FE_OFN34_write),
	.A(n96), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U13 (
	.ZN(n96),
	.A2(write),
	.A1(data[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U14 (
	.ZN(n63),
	.B2(n79),
	.B1(FE_OFN34_write),
	.A(n95), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U15 (
	.ZN(n95),
	.A2(FE_OFN34_write),
	.A1(data[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U16 (
	.ZN(n62),
	.B2(n78),
	.B1(write),
	.A(n94), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U17 (
	.ZN(n94),
	.A2(write),
	.A1(data[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U18 (
	.ZN(n61),
	.B2(n77),
	.B1(FE_OFN6_write),
	.A(n93), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U19 (
	.ZN(n93),
	.A2(FE_OFN6_write),
	.A1(data[8]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U20 (
	.ZN(n60),
	.B2(n76),
	.B1(FE_OFN34_write),
	.A(n92), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U21 (
	.ZN(n92),
	.A2(FE_OFN34_write),
	.A1(data[9]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U22 (
	.ZN(n59),
	.B2(n75),
	.B1(FE_OFN34_write),
	.A(n91), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U23 (
	.ZN(n91),
	.A2(FE_OFN34_write),
	.A1(data[10]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U24 (
	.ZN(n58),
	.B2(n74),
	.B1(FE_OFN34_write),
	.A(n90), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U25 (
	.ZN(n90),
	.A2(FE_OFN34_write),
	.A1(data[11]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U26 (
	.ZN(n57),
	.B2(n73),
	.B1(FE_OFN34_write),
	.A(n89), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U27 (
	.ZN(n89),
	.A2(FE_OFN34_write),
	.A1(data[12]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U28 (
	.ZN(n56),
	.B2(n72),
	.B1(FE_OFN6_write),
	.A(n88), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U29 (
	.ZN(n88),
	.A2(FE_OFN6_write),
	.A1(data[13]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U30 (
	.ZN(n55),
	.B2(n71),
	.B1(FE_OFN6_write),
	.A(n87), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U31 (
	.ZN(n87),
	.A2(FE_OFN6_write),
	.A1(data[14]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X2 U32 (
	.ZN(n54),
	.A(reset), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U33 (
	.ZN(n53),
	.B2(n70),
	.B1(FE_OFN6_write),
	.A(n86), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U34 (
	.ZN(n86),
	.A2(FE_OFN6_write),
	.A1(data[15]), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module SingleReg_21 (
	data, 
	clk, 
	reset, 
	write, 
	dataOut, 
	FE_OFN6_write, 
	FE_OFN7_write, 
	FE_OFN9_write, 
	FE_OFN40_write, 
	FE_OFN43_write, 
	FE_OFN45_write, 
	FE_OFN50_write, 
	clk__L2_N12, 
	VDD, 
	VSS);
   input [15:0] data;
   input clk;
   input reset;
   input write;
   output [15:0] dataOut;
   input FE_OFN6_write;
   input FE_OFN7_write;
   input FE_OFN9_write;
   input FE_OFN40_write;
   input FE_OFN43_write;
   input FE_OFN45_write;
   input FE_OFN50_write;
   input clk__L2_N12;
   inout VDD;
   inout VSS;

   // Internal wires
   wire n53;
   wire n54;
   wire n55;
   wire n56;
   wire n57;
   wire n58;
   wire n59;
   wire n60;
   wire n61;
   wire n62;
   wire n63;
   wire n64;
   wire n65;
   wire n66;
   wire n67;
   wire n68;
   wire n69;
   wire n70;
   wire n71;
   wire n72;
   wire n73;
   wire n74;
   wire n75;
   wire n76;
   wire n77;
   wire n78;
   wire n79;
   wire n80;
   wire n81;
   wire n82;
   wire n83;
   wire n84;
   wire n85;
   wire n86;
   wire n87;
   wire n88;
   wire n89;
   wire n90;
   wire n91;
   wire n92;
   wire n93;
   wire n94;
   wire n95;
   wire n96;
   wire n97;
   wire n98;
   wire n99;
   wire n100;
   wire n101;

   // Module instantiations
   DFFR_X1 \Reg_reg[15]  (
	.RN(n54),
	.QN(n70),
	.Q(dataOut[15]),
	.D(n53),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[14]  (
	.RN(n54),
	.QN(n71),
	.Q(dataOut[14]),
	.D(n55),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[13]  (
	.RN(n54),
	.QN(n72),
	.Q(dataOut[13]),
	.D(n56),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[12]  (
	.RN(n54),
	.QN(n73),
	.Q(dataOut[12]),
	.D(n57),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[11]  (
	.RN(n54),
	.QN(n74),
	.Q(dataOut[11]),
	.D(n58),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[10]  (
	.RN(n54),
	.QN(n75),
	.Q(dataOut[10]),
	.D(n59),
	.CK(clk__L2_N12), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[9]  (
	.RN(n54),
	.QN(n76),
	.Q(dataOut[9]),
	.D(n60),
	.CK(clk__L2_N12), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[8]  (
	.RN(n54),
	.QN(n77),
	.Q(dataOut[8]),
	.D(n61),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[7]  (
	.RN(n54),
	.QN(n78),
	.Q(dataOut[7]),
	.D(n62),
	.CK(clk__L2_N12), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[6]  (
	.RN(n54),
	.QN(n79),
	.Q(dataOut[6]),
	.D(n63),
	.CK(clk__L2_N12), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[5]  (
	.RN(n54),
	.QN(n80),
	.Q(dataOut[5]),
	.D(n64),
	.CK(clk__L2_N12), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[4]  (
	.RN(n54),
	.QN(n81),
	.Q(dataOut[4]),
	.D(n65),
	.CK(clk__L2_N12), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[3]  (
	.RN(n54),
	.QN(n82),
	.Q(dataOut[3]),
	.D(n66),
	.CK(clk__L2_N12), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[2]  (
	.RN(n54),
	.QN(n83),
	.Q(dataOut[2]),
	.D(n67),
	.CK(clk__L2_N12), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[1]  (
	.RN(n54),
	.QN(n84),
	.Q(dataOut[1]),
	.D(n68),
	.CK(clk__L2_N12), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[0]  (
	.RN(n54),
	.QN(n85),
	.Q(dataOut[0]),
	.D(n69),
	.CK(clk__L2_N12), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U2 (
	.ZN(n69),
	.B2(n85),
	.B1(FE_OFN40_write),
	.A(n101), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U3 (
	.ZN(n101),
	.A2(data[0]),
	.A1(FE_OFN43_write), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U4 (
	.ZN(n68),
	.B2(n84),
	.B1(FE_OFN40_write),
	.A(n100), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U5 (
	.ZN(n100),
	.A2(FE_OFN40_write),
	.A1(data[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U6 (
	.ZN(n67),
	.B2(n83),
	.B1(write),
	.A(n99), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U7 (
	.ZN(n99),
	.A2(write),
	.A1(data[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U8 (
	.ZN(n66),
	.B2(n82),
	.B1(FE_OFN40_write),
	.A(n98), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U9 (
	.ZN(n98),
	.A2(FE_OFN40_write),
	.A1(data[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U10 (
	.ZN(n65),
	.B2(n81),
	.B1(write),
	.A(n97), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U11 (
	.ZN(n97),
	.A2(FE_OFN9_write),
	.A1(data[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U12 (
	.ZN(n64),
	.B2(n80),
	.B1(write),
	.A(n96), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U13 (
	.ZN(n96),
	.A2(write),
	.A1(data[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U14 (
	.ZN(n63),
	.B2(n79),
	.B1(FE_OFN7_write),
	.A(n95), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U15 (
	.ZN(n95),
	.A2(FE_OFN7_write),
	.A1(data[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U16 (
	.ZN(n62),
	.B2(n78),
	.B1(write),
	.A(n94), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U17 (
	.ZN(n94),
	.A2(write),
	.A1(data[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U18 (
	.ZN(n61),
	.B2(n77),
	.B1(FE_OFN6_write),
	.A(n93), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U19 (
	.ZN(n93),
	.A2(FE_OFN6_write),
	.A1(data[8]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U20 (
	.ZN(n60),
	.B2(n76),
	.B1(FE_OFN7_write),
	.A(n92), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U21 (
	.ZN(n92),
	.A2(FE_OFN7_write),
	.A1(data[9]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U22 (
	.ZN(n59),
	.B2(n75),
	.B1(FE_OFN50_write),
	.A(n91), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U23 (
	.ZN(n91),
	.A2(FE_OFN50_write),
	.A1(data[10]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U24 (
	.ZN(n58),
	.B2(n74),
	.B1(FE_OFN7_write),
	.A(n90), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U25 (
	.ZN(n90),
	.A2(FE_OFN7_write),
	.A1(data[11]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U26 (
	.ZN(n57),
	.B2(n73),
	.B1(FE_OFN7_write),
	.A(n89), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U27 (
	.ZN(n89),
	.A2(FE_OFN7_write),
	.A1(data[12]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U28 (
	.ZN(n56),
	.B2(n72),
	.B1(FE_OFN45_write),
	.A(n88), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U29 (
	.ZN(n88),
	.A2(FE_OFN45_write),
	.A1(data[13]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U30 (
	.ZN(n55),
	.B2(n71),
	.B1(FE_OFN6_write),
	.A(n87), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U31 (
	.ZN(n87),
	.A2(FE_OFN6_write),
	.A1(data[14]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U32 (
	.ZN(n54),
	.A(reset), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U33 (
	.ZN(n53),
	.B2(n70),
	.B1(FE_OFN7_write),
	.A(n86), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U34 (
	.ZN(n86),
	.A2(FE_OFN7_write),
	.A1(data[15]), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module SingleReg_20 (
	data, 
	clk, 
	reset, 
	write, 
	dataOut, 
	FE_OFN6_write, 
	FE_OFN7_write, 
	FE_OFN34_write, 
	FE_OFN38_write, 
	FE_OFN40_write, 
	FE_OFN43_write, 
	FE_OFN45_write, 
	clk__L2_N12, 
	clk__L2_N2, 
	clk__L2_N6, 
	VDD, 
	VSS);
   input [15:0] data;
   input clk;
   input reset;
   input write;
   output [15:0] dataOut;
   input FE_OFN6_write;
   input FE_OFN7_write;
   input FE_OFN34_write;
   input FE_OFN38_write;
   input FE_OFN40_write;
   input FE_OFN43_write;
   input FE_OFN45_write;
   input clk__L2_N12;
   input clk__L2_N2;
   input clk__L2_N6;
   inout VDD;
   inout VSS;

   // Internal wires
   wire n53;
   wire n54;
   wire n55;
   wire n56;
   wire n57;
   wire n58;
   wire n59;
   wire n60;
   wire n61;
   wire n62;
   wire n63;
   wire n64;
   wire n65;
   wire n66;
   wire n67;
   wire n68;
   wire n69;
   wire n70;
   wire n71;
   wire n72;
   wire n73;
   wire n74;
   wire n75;
   wire n76;
   wire n77;
   wire n78;
   wire n79;
   wire n80;
   wire n81;
   wire n82;
   wire n83;
   wire n84;
   wire n85;
   wire n86;
   wire n87;
   wire n88;
   wire n89;
   wire n90;
   wire n91;
   wire n92;
   wire n93;
   wire n94;
   wire n95;
   wire n96;
   wire n97;
   wire n98;
   wire n99;
   wire n100;
   wire n101;

   // Module instantiations
   DFFR_X1 \Reg_reg[15]  (
	.RN(n54),
	.QN(n70),
	.Q(dataOut[15]),
	.D(n53),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[14]  (
	.RN(n54),
	.QN(n71),
	.Q(dataOut[14]),
	.D(n55),
	.CK(clk__L2_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[13]  (
	.RN(n54),
	.QN(n72),
	.Q(dataOut[13]),
	.D(n56),
	.CK(clk__L2_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[12]  (
	.RN(n54),
	.QN(n73),
	.Q(dataOut[12]),
	.D(n57),
	.CK(clk__L2_N12), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[11]  (
	.RN(n54),
	.QN(n74),
	.Q(dataOut[11]),
	.D(n58),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[10]  (
	.RN(n54),
	.QN(n75),
	.Q(dataOut[10]),
	.D(n59),
	.CK(clk__L2_N12), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[9]  (
	.RN(n54),
	.QN(n76),
	.Q(dataOut[9]),
	.D(n60),
	.CK(clk__L2_N12), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[8]  (
	.RN(n54),
	.QN(n77),
	.Q(dataOut[8]),
	.D(n61),
	.CK(clk__L2_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[7]  (
	.RN(n54),
	.QN(n78),
	.Q(dataOut[7]),
	.D(n62),
	.CK(clk__L2_N12), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[6]  (
	.RN(n54),
	.QN(n79),
	.Q(dataOut[6]),
	.D(n63),
	.CK(clk__L2_N12), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[5]  (
	.RN(n54),
	.QN(n80),
	.Q(dataOut[5]),
	.D(n64),
	.CK(clk__L2_N12), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[4]  (
	.RN(n54),
	.QN(n81),
	.Q(dataOut[4]),
	.D(n65),
	.CK(clk__L2_N12), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[3]  (
	.RN(n54),
	.QN(n82),
	.Q(dataOut[3]),
	.D(n66),
	.CK(clk__L2_N12), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[2]  (
	.RN(n54),
	.QN(n83),
	.Q(dataOut[2]),
	.D(n67),
	.CK(clk__L2_N12), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[1]  (
	.RN(n54),
	.QN(n84),
	.Q(dataOut[1]),
	.D(n68),
	.CK(clk__L2_N6), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[0]  (
	.RN(n54),
	.QN(n85),
	.Q(dataOut[0]),
	.D(n69),
	.CK(clk__L2_N6), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U2 (
	.ZN(n69),
	.B2(n85),
	.B1(FE_OFN40_write),
	.A(n101), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U3 (
	.ZN(n101),
	.A2(data[0]),
	.A1(FE_OFN40_write), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U4 (
	.ZN(n68),
	.B2(n84),
	.B1(FE_OFN40_write),
	.A(n100), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U5 (
	.ZN(n100),
	.A2(FE_OFN40_write),
	.A1(data[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U6 (
	.ZN(n67),
	.B2(n83),
	.B1(FE_OFN43_write),
	.A(n99), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U7 (
	.ZN(n99),
	.A2(FE_OFN43_write),
	.A1(data[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U8 (
	.ZN(n66),
	.B2(n82),
	.B1(FE_OFN43_write),
	.A(n98), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U9 (
	.ZN(n98),
	.A2(FE_OFN43_write),
	.A1(data[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U10 (
	.ZN(n65),
	.B2(n81),
	.B1(write),
	.A(n97), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U11 (
	.ZN(n97),
	.A2(write),
	.A1(data[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U12 (
	.ZN(n64),
	.B2(n80),
	.B1(write),
	.A(n96), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U13 (
	.ZN(n96),
	.A2(write),
	.A1(data[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U14 (
	.ZN(n63),
	.B2(n79),
	.B1(FE_OFN7_write),
	.A(n95), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U15 (
	.ZN(n95),
	.A2(FE_OFN38_write),
	.A1(data[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U16 (
	.ZN(n62),
	.B2(n78),
	.B1(write),
	.A(n94), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U17 (
	.ZN(n94),
	.A2(write),
	.A1(data[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U18 (
	.ZN(n61),
	.B2(n77),
	.B1(FE_OFN6_write),
	.A(n93), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U19 (
	.ZN(n93),
	.A2(FE_OFN6_write),
	.A1(data[8]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U20 (
	.ZN(n60),
	.B2(n76),
	.B1(FE_OFN38_write),
	.A(n92), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U21 (
	.ZN(n92),
	.A2(FE_OFN38_write),
	.A1(data[9]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U22 (
	.ZN(n59),
	.B2(n75),
	.B1(FE_OFN34_write),
	.A(n91), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U23 (
	.ZN(n91),
	.A2(FE_OFN34_write),
	.A1(data[10]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U24 (
	.ZN(n58),
	.B2(n74),
	.B1(FE_OFN7_write),
	.A(n90), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U25 (
	.ZN(n90),
	.A2(FE_OFN7_write),
	.A1(data[11]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U26 (
	.ZN(n57),
	.B2(n73),
	.B1(FE_OFN45_write),
	.A(n89), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U27 (
	.ZN(n89),
	.A2(FE_OFN45_write),
	.A1(data[12]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U28 (
	.ZN(n56),
	.B2(n72),
	.B1(FE_OFN6_write),
	.A(n88), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U29 (
	.ZN(n88),
	.A2(FE_OFN6_write),
	.A1(data[13]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U30 (
	.ZN(n55),
	.B2(n71),
	.B1(FE_OFN6_write),
	.A(n87), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U31 (
	.ZN(n87),
	.A2(FE_OFN6_write),
	.A1(data[14]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U32 (
	.ZN(n54),
	.A(reset), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U33 (
	.ZN(n53),
	.B2(n70),
	.B1(FE_OFN6_write),
	.A(n86), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U34 (
	.ZN(n86),
	.A2(FE_OFN6_write),
	.A1(data[15]), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module SingleReg_19 (
	data, 
	clk, 
	reset, 
	write, 
	dataOut, 
	FE_OFN7_write, 
	FE_OFN9_write, 
	FE_OFN50_write, 
	FE_OFN55_write, 
	clk__L2_N11, 
	clk__L2_N12, 
	clk__L2_N6, 
	VDD, 
	VSS);
   input [15:0] data;
   input clk;
   input reset;
   input write;
   output [15:0] dataOut;
   input FE_OFN7_write;
   input FE_OFN9_write;
   input FE_OFN50_write;
   input FE_OFN55_write;
   input clk__L2_N11;
   input clk__L2_N12;
   input clk__L2_N6;
   inout VDD;
   inout VSS;

   // Internal wires
   wire n53;
   wire n54;
   wire n55;
   wire n56;
   wire n57;
   wire n58;
   wire n59;
   wire n60;
   wire n61;
   wire n62;
   wire n63;
   wire n64;
   wire n65;
   wire n66;
   wire n67;
   wire n68;
   wire n69;
   wire n70;
   wire n71;
   wire n72;
   wire n73;
   wire n74;
   wire n75;
   wire n76;
   wire n77;
   wire n78;
   wire n79;
   wire n80;
   wire n81;
   wire n82;
   wire n83;
   wire n84;
   wire n85;
   wire n86;
   wire n87;
   wire n88;
   wire n89;
   wire n90;
   wire n91;
   wire n92;
   wire n93;
   wire n94;
   wire n95;
   wire n96;
   wire n97;
   wire n98;
   wire n99;
   wire n100;
   wire n101;

   // Module instantiations
   DFFR_X1 \Reg_reg[15]  (
	.RN(n54),
	.QN(n70),
	.Q(dataOut[15]),
	.D(n53),
	.CK(clk__L2_N11), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[14]  (
	.RN(n54),
	.QN(n71),
	.Q(dataOut[14]),
	.D(n55),
	.CK(clk__L2_N11), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[13]  (
	.RN(n54),
	.QN(n72),
	.Q(dataOut[13]),
	.D(n56),
	.CK(clk__L2_N11), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[12]  (
	.RN(n54),
	.QN(n73),
	.Q(dataOut[12]),
	.D(n57),
	.CK(clk__L2_N11), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[11]  (
	.RN(n54),
	.QN(n74),
	.Q(dataOut[11]),
	.D(n58),
	.CK(clk__L2_N11), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[10]  (
	.RN(n54),
	.QN(n75),
	.Q(dataOut[10]),
	.D(n59),
	.CK(clk__L2_N11), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[9]  (
	.RN(n54),
	.QN(n76),
	.Q(dataOut[9]),
	.D(n60),
	.CK(clk__L2_N12), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[8]  (
	.RN(n54),
	.QN(n77),
	.Q(dataOut[8]),
	.D(n61),
	.CK(clk__L2_N11), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[7]  (
	.RN(n54),
	.QN(n78),
	.Q(dataOut[7]),
	.D(n62),
	.CK(clk__L2_N11), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[6]  (
	.RN(n54),
	.QN(n79),
	.Q(dataOut[6]),
	.D(n63),
	.CK(clk__L2_N12), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[5]  (
	.RN(n54),
	.QN(n80),
	.Q(dataOut[5]),
	.D(n64),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[4]  (
	.RN(n54),
	.QN(n81),
	.Q(dataOut[4]),
	.D(n65),
	.CK(clk__L2_N12), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[3]  (
	.RN(n54),
	.QN(n82),
	.Q(dataOut[3]),
	.D(n66),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[2]  (
	.RN(n54),
	.QN(n83),
	.Q(dataOut[2]),
	.D(n67),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[1]  (
	.RN(n54),
	.QN(n84),
	.Q(dataOut[1]),
	.D(n68),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[0]  (
	.RN(n54),
	.QN(n85),
	.Q(dataOut[0]),
	.D(n69),
	.CK(clk__L2_N6), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U2 (
	.ZN(n69),
	.B2(n85),
	.B1(FE_OFN55_write),
	.A(n101), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U3 (
	.ZN(n101),
	.A2(data[0]),
	.A1(FE_OFN55_write), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U4 (
	.ZN(n68),
	.B2(n84),
	.B1(FE_OFN55_write),
	.A(n100), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U5 (
	.ZN(n100),
	.A2(FE_OFN55_write),
	.A1(data[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U6 (
	.ZN(n67),
	.B2(n83),
	.B1(FE_OFN55_write),
	.A(n99), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U7 (
	.ZN(n99),
	.A2(FE_OFN55_write),
	.A1(data[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U8 (
	.ZN(n66),
	.B2(n82),
	.B1(FE_OFN55_write),
	.A(n98), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U9 (
	.ZN(n98),
	.A2(FE_OFN55_write),
	.A1(data[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U10 (
	.ZN(n65),
	.B2(n81),
	.B1(FE_OFN55_write),
	.A(n97), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U11 (
	.ZN(n97),
	.A2(FE_OFN55_write),
	.A1(data[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U12 (
	.ZN(n64),
	.B2(n80),
	.B1(FE_OFN55_write),
	.A(n96), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U13 (
	.ZN(n96),
	.A2(FE_OFN55_write),
	.A1(data[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U14 (
	.ZN(n63),
	.B2(n79),
	.B1(FE_OFN7_write),
	.A(n95), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U15 (
	.ZN(n95),
	.A2(FE_OFN50_write),
	.A1(data[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U16 (
	.ZN(n62),
	.B2(n78),
	.B1(FE_OFN9_write),
	.A(n94), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U17 (
	.ZN(n94),
	.A2(FE_OFN50_write),
	.A1(data[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U18 (
	.ZN(n61),
	.B2(n77),
	.B1(write),
	.A(n93), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U19 (
	.ZN(n93),
	.A2(write),
	.A1(data[8]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U20 (
	.ZN(n60),
	.B2(n76),
	.B1(FE_OFN55_write),
	.A(n92), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U21 (
	.ZN(n92),
	.A2(FE_OFN55_write),
	.A1(data[9]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U22 (
	.ZN(n59),
	.B2(n75),
	.B1(FE_OFN50_write),
	.A(n91), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U23 (
	.ZN(n91),
	.A2(FE_OFN50_write),
	.A1(data[10]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U24 (
	.ZN(n58),
	.B2(n74),
	.B1(FE_OFN7_write),
	.A(n90), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U25 (
	.ZN(n90),
	.A2(FE_OFN7_write),
	.A1(data[11]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U26 (
	.ZN(n57),
	.B2(n73),
	.B1(FE_OFN7_write),
	.A(n89), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U27 (
	.ZN(n89),
	.A2(FE_OFN7_write),
	.A1(data[12]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U28 (
	.ZN(n56),
	.B2(n72),
	.B1(write),
	.A(n88), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U29 (
	.ZN(n88),
	.A2(write),
	.A1(data[13]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U30 (
	.ZN(n55),
	.B2(n71),
	.B1(write),
	.A(n87), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U31 (
	.ZN(n87),
	.A2(write),
	.A1(data[14]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X2 U32 (
	.ZN(n54),
	.A(reset), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U33 (
	.ZN(n53),
	.B2(n70),
	.B1(write),
	.A(n86), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U34 (
	.ZN(n86),
	.A2(write),
	.A1(data[15]), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module SingleReg_18 (
	data, 
	clk, 
	reset, 
	write, 
	dataOut, 
	FE_OFN7_write, 
	FE_OFN9_write, 
	FE_OFN50_write, 
	clk__L2_N11, 
	clk__L2_N12, 
	VDD, 
	VSS);
   input [15:0] data;
   input clk;
   input reset;
   input write;
   output [15:0] dataOut;
   input FE_OFN7_write;
   input FE_OFN9_write;
   input FE_OFN50_write;
   input clk__L2_N11;
   input clk__L2_N12;
   inout VDD;
   inout VSS;

   // Internal wires
   wire n53;
   wire n54;
   wire n55;
   wire n56;
   wire n57;
   wire n58;
   wire n59;
   wire n60;
   wire n61;
   wire n62;
   wire n63;
   wire n64;
   wire n65;
   wire n66;
   wire n67;
   wire n68;
   wire n69;
   wire n70;
   wire n71;
   wire n72;
   wire n73;
   wire n74;
   wire n75;
   wire n76;
   wire n77;
   wire n78;
   wire n79;
   wire n80;
   wire n81;
   wire n82;
   wire n83;
   wire n84;
   wire n85;
   wire n86;
   wire n87;
   wire n88;
   wire n89;
   wire n90;
   wire n91;
   wire n92;
   wire n93;
   wire n94;
   wire n95;
   wire n96;
   wire n97;
   wire n98;
   wire n99;
   wire n100;
   wire n101;

   // Module instantiations
   DFFR_X1 \Reg_reg[15]  (
	.RN(n54),
	.QN(n70),
	.Q(dataOut[15]),
	.D(n53),
	.CK(clk__L2_N11), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[14]  (
	.RN(n54),
	.QN(n71),
	.Q(dataOut[14]),
	.D(n55),
	.CK(clk__L2_N11), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[13]  (
	.RN(n54),
	.QN(n72),
	.Q(dataOut[13]),
	.D(n56),
	.CK(clk__L2_N11), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[12]  (
	.RN(n54),
	.QN(n73),
	.Q(dataOut[12]),
	.D(n57),
	.CK(clk__L2_N11), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[11]  (
	.RN(n54),
	.QN(n74),
	.Q(dataOut[11]),
	.D(n58),
	.CK(clk__L2_N11), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[10]  (
	.RN(n54),
	.QN(n75),
	.Q(dataOut[10]),
	.D(n59),
	.CK(clk__L2_N12), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[9]  (
	.RN(n54),
	.QN(n76),
	.Q(dataOut[9]),
	.D(n60),
	.CK(clk__L2_N12), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[8]  (
	.RN(n54),
	.QN(n77),
	.Q(dataOut[8]),
	.D(n61),
	.CK(clk__L2_N11), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[7]  (
	.RN(n54),
	.QN(n78),
	.Q(dataOut[7]),
	.D(n62),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[6]  (
	.RN(n54),
	.QN(n79),
	.Q(dataOut[6]),
	.D(n63),
	.CK(clk__L2_N12), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[5]  (
	.RN(n54),
	.QN(n80),
	.Q(dataOut[5]),
	.D(n64),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[4]  (
	.RN(n54),
	.QN(n81),
	.Q(dataOut[4]),
	.D(n65),
	.CK(clk__L2_N12), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[3]  (
	.RN(n54),
	.QN(n82),
	.Q(dataOut[3]),
	.D(n66),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[2]  (
	.RN(n54),
	.QN(n83),
	.Q(dataOut[2]),
	.D(n67),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[1]  (
	.RN(n54),
	.QN(n84),
	.Q(dataOut[1]),
	.D(n68),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[0]  (
	.RN(n54),
	.QN(n85),
	.Q(dataOut[0]),
	.D(n69),
	.CK(clk__L2_N12), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U2 (
	.ZN(n69),
	.B2(n85),
	.B1(FE_OFN9_write),
	.A(n101), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U3 (
	.ZN(n101),
	.A2(data[0]),
	.A1(FE_OFN9_write), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U4 (
	.ZN(n68),
	.B2(n84),
	.B1(FE_OFN9_write),
	.A(n100), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U5 (
	.ZN(n100),
	.A2(FE_OFN9_write),
	.A1(data[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U6 (
	.ZN(n67),
	.B2(n83),
	.B1(FE_OFN9_write),
	.A(n99), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U7 (
	.ZN(n99),
	.A2(FE_OFN9_write),
	.A1(data[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U8 (
	.ZN(n66),
	.B2(n82),
	.B1(FE_OFN9_write),
	.A(n98), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U9 (
	.ZN(n98),
	.A2(FE_OFN9_write),
	.A1(data[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U10 (
	.ZN(n65),
	.B2(n81),
	.B1(FE_OFN9_write),
	.A(n97), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U11 (
	.ZN(n97),
	.A2(FE_OFN9_write),
	.A1(data[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U12 (
	.ZN(n64),
	.B2(n80),
	.B1(FE_OFN9_write),
	.A(n96), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U13 (
	.ZN(n96),
	.A2(FE_OFN9_write),
	.A1(data[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U14 (
	.ZN(n63),
	.B2(n79),
	.B1(FE_OFN50_write),
	.A(n95), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U15 (
	.ZN(n95),
	.A2(FE_OFN50_write),
	.A1(data[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U16 (
	.ZN(n62),
	.B2(n78),
	.B1(FE_OFN9_write),
	.A(n94), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U17 (
	.ZN(n94),
	.A2(FE_OFN9_write),
	.A1(data[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U18 (
	.ZN(n61),
	.B2(n77),
	.B1(write),
	.A(n93), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U19 (
	.ZN(n93),
	.A2(write),
	.A1(data[8]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U20 (
	.ZN(n60),
	.B2(n76),
	.B1(FE_OFN9_write),
	.A(n92), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U21 (
	.ZN(n92),
	.A2(FE_OFN50_write),
	.A1(data[9]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U22 (
	.ZN(n59),
	.B2(n75),
	.B1(FE_OFN7_write),
	.A(n91), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U23 (
	.ZN(n91),
	.A2(FE_OFN7_write),
	.A1(data[10]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U24 (
	.ZN(n58),
	.B2(n74),
	.B1(FE_OFN7_write),
	.A(n90), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U25 (
	.ZN(n90),
	.A2(FE_OFN7_write),
	.A1(data[11]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U26 (
	.ZN(n57),
	.B2(n73),
	.B1(FE_OFN7_write),
	.A(n89), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U27 (
	.ZN(n89),
	.A2(FE_OFN7_write),
	.A1(data[12]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U28 (
	.ZN(n56),
	.B2(n72),
	.B1(write),
	.A(n88), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U29 (
	.ZN(n88),
	.A2(write),
	.A1(data[13]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U30 (
	.ZN(n55),
	.B2(n71),
	.B1(write),
	.A(n87), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U31 (
	.ZN(n87),
	.A2(FE_OFN7_write),
	.A1(data[14]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U32 (
	.ZN(n54),
	.A(reset), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U33 (
	.ZN(n53),
	.B2(n70),
	.B1(FE_OFN7_write),
	.A(n86), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U34 (
	.ZN(n86),
	.A2(FE_OFN7_write),
	.A1(data[15]), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module SingleReg_17 (
	data, 
	clk, 
	reset, 
	write, 
	dataOut, 
	FE_OFN9_write, 
	clk__L2_N11, 
	VDD, 
	VSS);
   input [15:0] data;
   input clk;
   input reset;
   input write;
   output [15:0] dataOut;
   input FE_OFN9_write;
   input clk__L2_N11;
   inout VDD;
   inout VSS;

   // Internal wires
   wire n53;
   wire n54;
   wire n55;
   wire n56;
   wire n57;
   wire n58;
   wire n59;
   wire n60;
   wire n61;
   wire n62;
   wire n63;
   wire n64;
   wire n65;
   wire n66;
   wire n67;
   wire n68;
   wire n69;
   wire n70;
   wire n71;
   wire n72;
   wire n73;
   wire n74;
   wire n75;
   wire n76;
   wire n77;
   wire n78;
   wire n79;
   wire n80;
   wire n81;
   wire n82;
   wire n83;
   wire n84;
   wire n85;
   wire n86;
   wire n87;
   wire n88;
   wire n89;
   wire n90;
   wire n91;
   wire n92;
   wire n93;
   wire n94;
   wire n95;
   wire n96;
   wire n97;
   wire n98;
   wire n99;
   wire n100;
   wire n101;

   // Module instantiations
   DFFR_X1 \Reg_reg[15]  (
	.RN(n54),
	.QN(n70),
	.Q(dataOut[15]),
	.D(n53),
	.CK(clk__L2_N11), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[14]  (
	.RN(n54),
	.QN(n71),
	.Q(dataOut[14]),
	.D(n55),
	.CK(clk__L2_N11), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[13]  (
	.RN(n54),
	.QN(n72),
	.Q(dataOut[13]),
	.D(n56),
	.CK(clk__L2_N11), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[12]  (
	.RN(n54),
	.QN(n73),
	.Q(dataOut[12]),
	.D(n57),
	.CK(clk__L2_N11), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[11]  (
	.RN(n54),
	.QN(n74),
	.Q(dataOut[11]),
	.D(n58),
	.CK(clk__L2_N11), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[10]  (
	.RN(n54),
	.QN(n75),
	.Q(dataOut[10]),
	.D(n59),
	.CK(clk__L2_N11), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[9]  (
	.RN(n54),
	.QN(n76),
	.Q(dataOut[9]),
	.D(n60),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[8]  (
	.RN(n54),
	.QN(n77),
	.Q(dataOut[8]),
	.D(n61),
	.CK(clk__L2_N11), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[7]  (
	.RN(n54),
	.QN(n78),
	.Q(dataOut[7]),
	.D(n62),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[6]  (
	.RN(n54),
	.QN(n79),
	.Q(dataOut[6]),
	.D(n63),
	.CK(clk__L2_N11), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[5]  (
	.RN(n54),
	.QN(n80),
	.Q(dataOut[5]),
	.D(n64),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[4]  (
	.RN(n54),
	.QN(n81),
	.Q(dataOut[4]),
	.D(n65),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[3]  (
	.RN(n54),
	.QN(n82),
	.Q(dataOut[3]),
	.D(n66),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[2]  (
	.RN(n54),
	.QN(n83),
	.Q(dataOut[2]),
	.D(n67),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[1]  (
	.RN(n54),
	.QN(n84),
	.Q(dataOut[1]),
	.D(n68),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[0]  (
	.RN(n54),
	.QN(n85),
	.Q(dataOut[0]),
	.D(n69),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U2 (
	.ZN(n69),
	.B2(n85),
	.B1(FE_OFN9_write),
	.A(n101), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U3 (
	.ZN(n101),
	.A2(data[0]),
	.A1(FE_OFN9_write), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U4 (
	.ZN(n68),
	.B2(n84),
	.B1(FE_OFN9_write),
	.A(n100), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U5 (
	.ZN(n100),
	.A2(FE_OFN9_write),
	.A1(data[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U6 (
	.ZN(n67),
	.B2(n83),
	.B1(FE_OFN9_write),
	.A(n99), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U7 (
	.ZN(n99),
	.A2(FE_OFN9_write),
	.A1(data[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U8 (
	.ZN(n66),
	.B2(n82),
	.B1(FE_OFN9_write),
	.A(n98), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U9 (
	.ZN(n98),
	.A2(FE_OFN9_write),
	.A1(data[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U10 (
	.ZN(n65),
	.B2(n81),
	.B1(FE_OFN9_write),
	.A(n97), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U11 (
	.ZN(n97),
	.A2(FE_OFN9_write),
	.A1(data[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U12 (
	.ZN(n64),
	.B2(n80),
	.B1(FE_OFN9_write),
	.A(n96), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U13 (
	.ZN(n96),
	.A2(FE_OFN9_write),
	.A1(data[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U14 (
	.ZN(n63),
	.B2(n79),
	.B1(write),
	.A(n95), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U15 (
	.ZN(n95),
	.A2(write),
	.A1(data[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U16 (
	.ZN(n62),
	.B2(n78),
	.B1(FE_OFN9_write),
	.A(n94), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U17 (
	.ZN(n94),
	.A2(FE_OFN9_write),
	.A1(data[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U18 (
	.ZN(n61),
	.B2(n77),
	.B1(write),
	.A(n93), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U19 (
	.ZN(n93),
	.A2(write),
	.A1(data[8]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U20 (
	.ZN(n60),
	.B2(n76),
	.B1(write),
	.A(n92), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U21 (
	.ZN(n92),
	.A2(write),
	.A1(data[9]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U22 (
	.ZN(n59),
	.B2(n75),
	.B1(write),
	.A(n91), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U23 (
	.ZN(n91),
	.A2(write),
	.A1(data[10]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U24 (
	.ZN(n58),
	.B2(n74),
	.B1(write),
	.A(n90), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U25 (
	.ZN(n90),
	.A2(write),
	.A1(data[11]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U26 (
	.ZN(n57),
	.B2(n73),
	.B1(write),
	.A(n89), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U27 (
	.ZN(n89),
	.A2(write),
	.A1(data[12]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U28 (
	.ZN(n56),
	.B2(n72),
	.B1(write),
	.A(n88), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U29 (
	.ZN(n88),
	.A2(write),
	.A1(data[13]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U30 (
	.ZN(n55),
	.B2(n71),
	.B1(write),
	.A(n87), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U31 (
	.ZN(n87),
	.A2(write),
	.A1(data[14]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U32 (
	.ZN(n54),
	.A(reset), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U33 (
	.ZN(n53),
	.B2(n70),
	.B1(write),
	.A(n86), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U34 (
	.ZN(n86),
	.A2(write),
	.A1(data[15]), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module SingleReg_16 (
	data, 
	clk, 
	reset, 
	write, 
	dataOut, 
	FE_OFN7_write, 
	FE_OFN9_write, 
	clk__L2_N11, 
	VDD, 
	VSS);
   input [15:0] data;
   input clk;
   input reset;
   input write;
   output [15:0] dataOut;
   input FE_OFN7_write;
   input FE_OFN9_write;
   input clk__L2_N11;
   inout VDD;
   inout VSS;

   // Internal wires
   wire FE_OFN52_write;
   wire n53;
   wire n54;
   wire n55;
   wire n56;
   wire n57;
   wire n58;
   wire n59;
   wire n60;
   wire n61;
   wire n62;
   wire n63;
   wire n64;
   wire n65;
   wire n66;
   wire n67;
   wire n68;
   wire n69;
   wire n70;
   wire n71;
   wire n72;
   wire n73;
   wire n74;
   wire n75;
   wire n76;
   wire n77;
   wire n78;
   wire n79;
   wire n80;
   wire n81;
   wire n82;
   wire n83;
   wire n84;
   wire n85;
   wire n86;
   wire n87;
   wire n88;
   wire n89;
   wire n90;
   wire n91;
   wire n92;
   wire n93;
   wire n94;
   wire n95;
   wire n96;
   wire n97;
   wire n98;
   wire n99;
   wire n100;
   wire n101;

   // Module instantiations
   BUF_X1 FE_OFC52_write (
	.Z(FE_OFN52_write),
	.A(FE_OFN7_write), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[15]  (
	.RN(n54),
	.QN(n70),
	.Q(dataOut[15]),
	.D(n53),
	.CK(clk__L2_N11), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[14]  (
	.RN(n54),
	.QN(n71),
	.Q(dataOut[14]),
	.D(n55),
	.CK(clk__L2_N11), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[13]  (
	.RN(n54),
	.QN(n72),
	.Q(dataOut[13]),
	.D(n56),
	.CK(clk__L2_N11), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[12]  (
	.RN(n54),
	.QN(n73),
	.Q(dataOut[12]),
	.D(n57),
	.CK(clk__L2_N11), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[11]  (
	.RN(n54),
	.QN(n74),
	.Q(dataOut[11]),
	.D(n58),
	.CK(clk__L2_N11), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[10]  (
	.RN(n54),
	.QN(n75),
	.Q(dataOut[10]),
	.D(n59),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[9]  (
	.RN(n54),
	.QN(n76),
	.Q(dataOut[9]),
	.D(n60),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[8]  (
	.RN(n54),
	.QN(n77),
	.Q(dataOut[8]),
	.D(n61),
	.CK(clk__L2_N11), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[7]  (
	.RN(n54),
	.QN(n78),
	.Q(dataOut[7]),
	.D(n62),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[6]  (
	.RN(n54),
	.QN(n79),
	.Q(dataOut[6]),
	.D(n63),
	.CK(clk__L2_N11), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[5]  (
	.RN(n54),
	.QN(n80),
	.Q(dataOut[5]),
	.D(n64),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[4]  (
	.RN(n54),
	.QN(n81),
	.Q(dataOut[4]),
	.D(n65),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[3]  (
	.RN(n54),
	.QN(n82),
	.Q(dataOut[3]),
	.D(n66),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[2]  (
	.RN(n54),
	.QN(n83),
	.Q(dataOut[2]),
	.D(n67),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[1]  (
	.RN(n54),
	.QN(n84),
	.Q(dataOut[1]),
	.D(n68),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[0]  (
	.RN(n54),
	.QN(n85),
	.Q(dataOut[0]),
	.D(n69),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U2 (
	.ZN(n69),
	.B2(n85),
	.B1(FE_OFN9_write),
	.A(n101), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U3 (
	.ZN(n101),
	.A2(data[0]),
	.A1(FE_OFN9_write), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U4 (
	.ZN(n68),
	.B2(n84),
	.B1(FE_OFN9_write),
	.A(n100), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U5 (
	.ZN(n100),
	.A2(FE_OFN9_write),
	.A1(data[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U6 (
	.ZN(n67),
	.B2(n83),
	.B1(FE_OFN9_write),
	.A(n99), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U7 (
	.ZN(n99),
	.A2(FE_OFN9_write),
	.A1(data[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U8 (
	.ZN(n66),
	.B2(n82),
	.B1(FE_OFN9_write),
	.A(n98), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U9 (
	.ZN(n98),
	.A2(FE_OFN9_write),
	.A1(data[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U10 (
	.ZN(n65),
	.B2(n81),
	.B1(FE_OFN9_write),
	.A(n97), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U11 (
	.ZN(n97),
	.A2(FE_OFN9_write),
	.A1(data[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U12 (
	.ZN(n64),
	.B2(n80),
	.B1(FE_OFN9_write),
	.A(n96), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U13 (
	.ZN(n96),
	.A2(FE_OFN9_write),
	.A1(data[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U14 (
	.ZN(n63),
	.B2(n79),
	.B1(FE_OFN7_write),
	.A(n95), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U15 (
	.ZN(n95),
	.A2(FE_OFN7_write),
	.A1(data[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U16 (
	.ZN(n62),
	.B2(n78),
	.B1(FE_OFN9_write),
	.A(n94), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U17 (
	.ZN(n94),
	.A2(FE_OFN9_write),
	.A1(data[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U18 (
	.ZN(n61),
	.B2(n77),
	.B1(FE_OFN52_write),
	.A(n93), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U19 (
	.ZN(n93),
	.A2(FE_OFN52_write),
	.A1(data[8]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U20 (
	.ZN(n60),
	.B2(n76),
	.B1(FE_OFN9_write),
	.A(n92), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U21 (
	.ZN(n92),
	.A2(FE_OFN9_write),
	.A1(data[9]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U22 (
	.ZN(n59),
	.B2(n75),
	.B1(FE_OFN7_write),
	.A(n91), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U23 (
	.ZN(n91),
	.A2(FE_OFN7_write),
	.A1(data[10]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U24 (
	.ZN(n58),
	.B2(n74),
	.B1(FE_OFN7_write),
	.A(n90), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U25 (
	.ZN(n90),
	.A2(FE_OFN7_write),
	.A1(data[11]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U26 (
	.ZN(n57),
	.B2(n73),
	.B1(FE_OFN7_write),
	.A(n89), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U27 (
	.ZN(n89),
	.A2(FE_OFN7_write),
	.A1(data[12]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U28 (
	.ZN(n56),
	.B2(n72),
	.B1(FE_OFN52_write),
	.A(n88), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U29 (
	.ZN(n88),
	.A2(FE_OFN52_write),
	.A1(data[13]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U30 (
	.ZN(n55),
	.B2(n71),
	.B1(write),
	.A(n87), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U31 (
	.ZN(n87),
	.A2(write),
	.A1(data[14]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U32 (
	.ZN(n54),
	.A(reset), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U33 (
	.ZN(n53),
	.B2(n70),
	.B1(FE_OFN7_write),
	.A(n86), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U34 (
	.ZN(n86),
	.A2(FE_OFN7_write),
	.A1(data[15]), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module SingleReg_15 (
	data, 
	clk, 
	reset, 
	write, 
	dataOut, 
	FE_OFN12_write, 
	FE_OFN3_write, 
	FE_OFN8_write, 
	FE_OFN26_write, 
	FE_OFN30_write, 
	clk__L2_N13, 
	clk__L2_N4, 
	clk__L2_N8, 
	VDD, 
	VSS);
   input [15:0] data;
   input clk;
   input reset;
   input write;
   output [15:0] dataOut;
   input FE_OFN12_write;
   input FE_OFN3_write;
   input FE_OFN8_write;
   input FE_OFN26_write;
   input FE_OFN30_write;
   input clk__L2_N13;
   input clk__L2_N4;
   input clk__L2_N8;
   inout VDD;
   inout VSS;

   // Internal wires
   wire n53;
   wire n54;
   wire n55;
   wire n56;
   wire n57;
   wire n58;
   wire n59;
   wire n60;
   wire n61;
   wire n62;
   wire n63;
   wire n64;
   wire n65;
   wire n66;
   wire n67;
   wire n68;
   wire n69;
   wire n70;
   wire n71;
   wire n72;
   wire n73;
   wire n74;
   wire n75;
   wire n76;
   wire n77;
   wire n78;
   wire n79;
   wire n80;
   wire n81;
   wire n82;
   wire n83;
   wire n84;
   wire n85;
   wire n86;
   wire n87;
   wire n88;
   wire n89;
   wire n90;
   wire n91;
   wire n92;
   wire n93;
   wire n94;
   wire n95;
   wire n96;
   wire n97;
   wire n98;
   wire n99;
   wire n100;
   wire n101;

   // Module instantiations
   DFFR_X1 \Reg_reg[15]  (
	.RN(n54),
	.QN(n70),
	.Q(dataOut[15]),
	.D(n53),
	.CK(clk__L2_N8), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[14]  (
	.RN(n54),
	.QN(n71),
	.Q(dataOut[14]),
	.D(n55),
	.CK(clk__L2_N8), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[13]  (
	.RN(n54),
	.QN(n72),
	.Q(dataOut[13]),
	.D(n56),
	.CK(clk__L2_N4), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[12]  (
	.RN(n54),
	.QN(n73),
	.Q(dataOut[12]),
	.D(n57),
	.CK(clk__L2_N8), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[11]  (
	.RN(n54),
	.QN(n74),
	.Q(dataOut[11]),
	.D(n58),
	.CK(clk__L2_N13), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[10]  (
	.RN(n54),
	.QN(n75),
	.Q(dataOut[10]),
	.D(n59),
	.CK(clk__L2_N4), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[9]  (
	.RN(n54),
	.QN(n76),
	.Q(dataOut[9]),
	.D(n60),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[8]  (
	.RN(n54),
	.QN(n77),
	.Q(dataOut[8]),
	.D(n61),
	.CK(clk__L2_N4), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[7]  (
	.RN(n54),
	.QN(n78),
	.Q(dataOut[7]),
	.D(n62),
	.CK(clk__L2_N13), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[6]  (
	.RN(n54),
	.QN(n79),
	.Q(dataOut[6]),
	.D(n63),
	.CK(clk__L2_N8), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[5]  (
	.RN(n54),
	.QN(n80),
	.Q(dataOut[5]),
	.D(n64),
	.CK(clk__L2_N13), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[4]  (
	.RN(n54),
	.QN(n81),
	.Q(dataOut[4]),
	.D(n65),
	.CK(clk__L2_N13), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[3]  (
	.RN(n54),
	.QN(n82),
	.Q(dataOut[3]),
	.D(n66),
	.CK(clk__L2_N13), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[2]  (
	.RN(n54),
	.QN(n83),
	.Q(dataOut[2]),
	.D(n67),
	.CK(clk__L2_N13), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[1]  (
	.RN(n54),
	.QN(n84),
	.Q(dataOut[1]),
	.D(n68),
	.CK(clk__L2_N13), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[0]  (
	.RN(n54),
	.QN(n85),
	.Q(dataOut[0]),
	.D(n69),
	.CK(clk__L2_N13), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U2 (
	.ZN(n69),
	.B2(n85),
	.B1(FE_OFN12_write),
	.A(n101), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U3 (
	.ZN(n101),
	.A2(data[0]),
	.A1(FE_OFN12_write), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U4 (
	.ZN(n68),
	.B2(n84),
	.B1(FE_OFN12_write),
	.A(n100), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U5 (
	.ZN(n100),
	.A2(FE_OFN12_write),
	.A1(data[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U6 (
	.ZN(n67),
	.B2(n83),
	.B1(FE_OFN12_write),
	.A(n99), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U7 (
	.ZN(n99),
	.A2(FE_OFN12_write),
	.A1(data[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U8 (
	.ZN(n66),
	.B2(n82),
	.B1(FE_OFN12_write),
	.A(n98), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U9 (
	.ZN(n98),
	.A2(FE_OFN12_write),
	.A1(data[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U10 (
	.ZN(n65),
	.B2(n81),
	.B1(FE_OFN26_write),
	.A(n97), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U11 (
	.ZN(n97),
	.A2(FE_OFN26_write),
	.A1(data[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U12 (
	.ZN(n64),
	.B2(n80),
	.B1(FE_OFN26_write),
	.A(n96), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U13 (
	.ZN(n96),
	.A2(FE_OFN26_write),
	.A1(data[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U14 (
	.ZN(n63),
	.B2(n79),
	.B1(FE_OFN26_write),
	.A(n95), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U15 (
	.ZN(n95),
	.A2(FE_OFN26_write),
	.A1(data[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U16 (
	.ZN(n62),
	.B2(n78),
	.B1(FE_OFN12_write),
	.A(n94), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U17 (
	.ZN(n94),
	.A2(FE_OFN12_write),
	.A1(data[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U18 (
	.ZN(n61),
	.B2(n77),
	.B1(FE_OFN8_write),
	.A(n93), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U19 (
	.ZN(n93),
	.A2(FE_OFN30_write),
	.A1(data[8]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U20 (
	.ZN(n60),
	.B2(n76),
	.B1(FE_OFN12_write),
	.A(n92), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U21 (
	.ZN(n92),
	.A2(FE_OFN12_write),
	.A1(data[9]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U22 (
	.ZN(n59),
	.B2(n75),
	.B1(FE_OFN8_write),
	.A(n91), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U23 (
	.ZN(n91),
	.A2(FE_OFN8_write),
	.A1(data[10]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U24 (
	.ZN(n58),
	.B2(n74),
	.B1(FE_OFN30_write),
	.A(n90), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U25 (
	.ZN(n90),
	.A2(FE_OFN30_write),
	.A1(data[11]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U26 (
	.ZN(n57),
	.B2(n73),
	.B1(FE_OFN3_write),
	.A(n89), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U27 (
	.ZN(n89),
	.A2(FE_OFN30_write),
	.A1(data[12]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U28 (
	.ZN(n56),
	.B2(n72),
	.B1(write),
	.A(n88), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U29 (
	.ZN(n88),
	.A2(write),
	.A1(data[13]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U30 (
	.ZN(n55),
	.B2(n71),
	.B1(write),
	.A(n87), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U31 (
	.ZN(n87),
	.A2(write),
	.A1(data[14]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X2 U32 (
	.ZN(n54),
	.A(reset), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U33 (
	.ZN(n53),
	.B2(n70),
	.B1(write),
	.A(n86), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U34 (
	.ZN(n86),
	.A2(write),
	.A1(data[15]), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module SingleReg_14 (
	data, 
	clk, 
	reset, 
	write, 
	dataOut, 
	FE_OFN10_write, 
	FE_OFN12_write, 
	FE_OFN3_write, 
	FE_OFN8_write, 
	FE_OFN30_write, 
	clk__L2_N4, 
	clk__L2_N8, 
	VDD, 
	VSS);
   input [15:0] data;
   input clk;
   input reset;
   input write;
   output [15:0] dataOut;
   input FE_OFN10_write;
   input FE_OFN12_write;
   input FE_OFN3_write;
   input FE_OFN8_write;
   input FE_OFN30_write;
   input clk__L2_N4;
   input clk__L2_N8;
   inout VDD;
   inout VSS;

   // Internal wires
   wire n53;
   wire n54;
   wire n55;
   wire n56;
   wire n57;
   wire n58;
   wire n59;
   wire n60;
   wire n61;
   wire n62;
   wire n63;
   wire n64;
   wire n65;
   wire n66;
   wire n67;
   wire n68;
   wire n69;
   wire n70;
   wire n71;
   wire n72;
   wire n73;
   wire n74;
   wire n75;
   wire n76;
   wire n77;
   wire n78;
   wire n79;
   wire n80;
   wire n81;
   wire n82;
   wire n83;
   wire n84;
   wire n85;
   wire n86;
   wire n87;
   wire n88;
   wire n89;
   wire n90;
   wire n91;
   wire n92;
   wire n93;
   wire n94;
   wire n95;
   wire n96;
   wire n97;
   wire n98;
   wire n99;
   wire n100;
   wire n101;

   // Module instantiations
   DFFR_X1 \Reg_reg[15]  (
	.RN(n54),
	.QN(n70),
	.Q(dataOut[15]),
	.D(n53),
	.CK(clk__L2_N8), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[14]  (
	.RN(n54),
	.QN(n71),
	.Q(dataOut[14]),
	.D(n55),
	.CK(clk__L2_N8), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[13]  (
	.RN(n54),
	.QN(n72),
	.Q(dataOut[13]),
	.D(n56),
	.CK(clk__L2_N4), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[12]  (
	.RN(n54),
	.QN(n73),
	.Q(dataOut[12]),
	.D(n57),
	.CK(clk__L2_N8), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[11]  (
	.RN(n54),
	.QN(n74),
	.Q(dataOut[11]),
	.D(n58),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[10]  (
	.RN(n54),
	.QN(n75),
	.Q(dataOut[10]),
	.D(n59),
	.CK(clk__L2_N4), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[9]  (
	.RN(n54),
	.QN(n76),
	.Q(dataOut[9]),
	.D(n60),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[8]  (
	.RN(n54),
	.QN(n77),
	.Q(dataOut[8]),
	.D(n61),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[7]  (
	.RN(n54),
	.QN(n78),
	.Q(dataOut[7]),
	.D(n62),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[6]  (
	.RN(n54),
	.QN(n79),
	.Q(dataOut[6]),
	.D(n63),
	.CK(clk__L2_N4), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[5]  (
	.RN(n54),
	.QN(n80),
	.Q(dataOut[5]),
	.D(n64),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[4]  (
	.RN(n54),
	.QN(n81),
	.Q(dataOut[4]),
	.D(n65),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[3]  (
	.RN(n54),
	.QN(n82),
	.Q(dataOut[3]),
	.D(n66),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[2]  (
	.RN(n54),
	.QN(n83),
	.Q(dataOut[2]),
	.D(n67),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[1]  (
	.RN(n54),
	.QN(n84),
	.Q(dataOut[1]),
	.D(n68),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[0]  (
	.RN(n54),
	.QN(n85),
	.Q(dataOut[0]),
	.D(n69),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U2 (
	.ZN(n69),
	.B2(n85),
	.B1(FE_OFN12_write),
	.A(n101), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U3 (
	.ZN(n101),
	.A2(data[0]),
	.A1(FE_OFN12_write), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U4 (
	.ZN(n68),
	.B2(n84),
	.B1(FE_OFN12_write),
	.A(n100), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U5 (
	.ZN(n100),
	.A2(FE_OFN12_write),
	.A1(data[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U6 (
	.ZN(n67),
	.B2(n83),
	.B1(FE_OFN12_write),
	.A(n99), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U7 (
	.ZN(n99),
	.A2(FE_OFN12_write),
	.A1(data[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U8 (
	.ZN(n66),
	.B2(n82),
	.B1(FE_OFN3_write),
	.A(n98), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U9 (
	.ZN(n98),
	.A2(FE_OFN3_write),
	.A1(data[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U10 (
	.ZN(n65),
	.B2(n81),
	.B1(FE_OFN3_write),
	.A(n97), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U11 (
	.ZN(n97),
	.A2(FE_OFN3_write),
	.A1(data[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U12 (
	.ZN(n64),
	.B2(n80),
	.B1(FE_OFN3_write),
	.A(n96), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U13 (
	.ZN(n96),
	.A2(FE_OFN3_write),
	.A1(data[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U14 (
	.ZN(n63),
	.B2(n79),
	.B1(FE_OFN3_write),
	.A(n95), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U15 (
	.ZN(n95),
	.A2(FE_OFN3_write),
	.A1(data[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U16 (
	.ZN(n62),
	.B2(n78),
	.B1(FE_OFN12_write),
	.A(n94), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U17 (
	.ZN(n94),
	.A2(FE_OFN12_write),
	.A1(data[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U18 (
	.ZN(n61),
	.B2(n77),
	.B1(FE_OFN30_write),
	.A(n93), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U19 (
	.ZN(n93),
	.A2(FE_OFN30_write),
	.A1(data[8]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U20 (
	.ZN(n60),
	.B2(n76),
	.B1(FE_OFN10_write),
	.A(n92), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U21 (
	.ZN(n92),
	.A2(FE_OFN10_write),
	.A1(data[9]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U22 (
	.ZN(n59),
	.B2(n75),
	.B1(FE_OFN8_write),
	.A(n91), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U23 (
	.ZN(n91),
	.A2(FE_OFN8_write),
	.A1(data[10]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U24 (
	.ZN(n58),
	.B2(n74),
	.B1(FE_OFN3_write),
	.A(n90), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U25 (
	.ZN(n90),
	.A2(FE_OFN30_write),
	.A1(data[11]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U26 (
	.ZN(n57),
	.B2(n73),
	.B1(FE_OFN30_write),
	.A(n89), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U27 (
	.ZN(n89),
	.A2(FE_OFN30_write),
	.A1(data[12]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U28 (
	.ZN(n56),
	.B2(n72),
	.B1(FE_OFN8_write),
	.A(n88), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U29 (
	.ZN(n88),
	.A2(FE_OFN8_write),
	.A1(data[13]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U30 (
	.ZN(n55),
	.B2(n71),
	.B1(FE_OFN8_write),
	.A(n87), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U31 (
	.ZN(n87),
	.A2(FE_OFN8_write),
	.A1(data[14]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U32 (
	.ZN(n54),
	.A(reset), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U33 (
	.ZN(n53),
	.B2(n70),
	.B1(write),
	.A(n86), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U34 (
	.ZN(n86),
	.A2(write),
	.A1(data[15]), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module SingleReg_13 (
	data, 
	clk, 
	reset, 
	write, 
	dataOut, 
	FE_OFN3_write, 
	FE_OFN28_write, 
	clk__L2_N8, 
	VDD, 
	VSS);
   input [15:0] data;
   input clk;
   input reset;
   input write;
   output [15:0] dataOut;
   input FE_OFN3_write;
   input FE_OFN28_write;
   input clk__L2_N8;
   inout VDD;
   inout VSS;

   // Internal wires
   wire n53;
   wire n54;
   wire n55;
   wire n56;
   wire n57;
   wire n58;
   wire n59;
   wire n60;
   wire n61;
   wire n62;
   wire n63;
   wire n64;
   wire n65;
   wire n66;
   wire n67;
   wire n68;
   wire n69;
   wire n70;
   wire n71;
   wire n72;
   wire n73;
   wire n74;
   wire n75;
   wire n76;
   wire n77;
   wire n78;
   wire n79;
   wire n80;
   wire n81;
   wire n82;
   wire n83;
   wire n84;
   wire n85;
   wire n86;
   wire n87;
   wire n88;
   wire n89;
   wire n90;
   wire n91;
   wire n92;
   wire n93;
   wire n94;
   wire n95;
   wire n96;
   wire n97;
   wire n98;
   wire n99;
   wire n100;
   wire n101;

   // Module instantiations
   DFFR_X1 \Reg_reg[15]  (
	.RN(n54),
	.QN(n70),
	.Q(dataOut[15]),
	.D(n53),
	.CK(clk__L2_N8), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[14]  (
	.RN(n54),
	.QN(n71),
	.Q(dataOut[14]),
	.D(n55),
	.CK(clk__L2_N8), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[13]  (
	.RN(n54),
	.QN(n72),
	.Q(dataOut[13]),
	.D(n56),
	.CK(clk__L2_N8), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[12]  (
	.RN(n54),
	.QN(n73),
	.Q(dataOut[12]),
	.D(n57),
	.CK(clk__L2_N8), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[11]  (
	.RN(n54),
	.QN(n74),
	.Q(dataOut[11]),
	.D(n58),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[10]  (
	.RN(n54),
	.QN(n75),
	.Q(dataOut[10]),
	.D(n59),
	.CK(clk__L2_N8), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[9]  (
	.RN(n54),
	.QN(n76),
	.Q(dataOut[9]),
	.D(n60),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[8]  (
	.RN(n54),
	.QN(n77),
	.Q(dataOut[8]),
	.D(n61),
	.CK(clk__L2_N8), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[7]  (
	.RN(n54),
	.QN(n78),
	.Q(dataOut[7]),
	.D(n62),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[6]  (
	.RN(n54),
	.QN(n79),
	.Q(dataOut[6]),
	.D(n63),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[5]  (
	.RN(n54),
	.QN(n80),
	.Q(dataOut[5]),
	.D(n64),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[4]  (
	.RN(n54),
	.QN(n81),
	.Q(dataOut[4]),
	.D(n65),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[3]  (
	.RN(n54),
	.QN(n82),
	.Q(dataOut[3]),
	.D(n66),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[2]  (
	.RN(n54),
	.QN(n83),
	.Q(dataOut[2]),
	.D(n67),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[1]  (
	.RN(n54),
	.QN(n84),
	.Q(dataOut[1]),
	.D(n68),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[0]  (
	.RN(n54),
	.QN(n85),
	.Q(dataOut[0]),
	.D(n69),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U2 (
	.ZN(n69),
	.B2(n85),
	.B1(FE_OFN28_write),
	.A(n101), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U3 (
	.ZN(n101),
	.A2(data[0]),
	.A1(FE_OFN28_write), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U4 (
	.ZN(n68),
	.B2(n84),
	.B1(FE_OFN28_write),
	.A(n100), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U5 (
	.ZN(n100),
	.A2(FE_OFN28_write),
	.A1(data[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U6 (
	.ZN(n67),
	.B2(n83),
	.B1(FE_OFN28_write),
	.A(n99), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U7 (
	.ZN(n99),
	.A2(FE_OFN28_write),
	.A1(data[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U8 (
	.ZN(n66),
	.B2(n82),
	.B1(FE_OFN28_write),
	.A(n98), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U9 (
	.ZN(n98),
	.A2(FE_OFN28_write),
	.A1(data[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U10 (
	.ZN(n65),
	.B2(n81),
	.B1(FE_OFN28_write),
	.A(n97), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U11 (
	.ZN(n97),
	.A2(FE_OFN28_write),
	.A1(data[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U12 (
	.ZN(n64),
	.B2(n80),
	.B1(FE_OFN28_write),
	.A(n96), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U13 (
	.ZN(n96),
	.A2(FE_OFN28_write),
	.A1(data[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U14 (
	.ZN(n63),
	.B2(n79),
	.B1(FE_OFN28_write),
	.A(n95), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U15 (
	.ZN(n95),
	.A2(FE_OFN28_write),
	.A1(data[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U16 (
	.ZN(n62),
	.B2(n78),
	.B1(FE_OFN28_write),
	.A(n94), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U17 (
	.ZN(n94),
	.A2(FE_OFN28_write),
	.A1(data[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U18 (
	.ZN(n61),
	.B2(n77),
	.B1(FE_OFN28_write),
	.A(n93), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U19 (
	.ZN(n93),
	.A2(FE_OFN28_write),
	.A1(data[8]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U20 (
	.ZN(n60),
	.B2(n76),
	.B1(FE_OFN28_write),
	.A(n92), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U21 (
	.ZN(n92),
	.A2(FE_OFN28_write),
	.A1(data[9]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U22 (
	.ZN(n59),
	.B2(n75),
	.B1(FE_OFN28_write),
	.A(n91), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U23 (
	.ZN(n91),
	.A2(FE_OFN28_write),
	.A1(data[10]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U24 (
	.ZN(n58),
	.B2(n74),
	.B1(FE_OFN3_write),
	.A(n90), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U25 (
	.ZN(n90),
	.A2(FE_OFN3_write),
	.A1(data[11]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U26 (
	.ZN(n57),
	.B2(n73),
	.B1(write),
	.A(n89), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U27 (
	.ZN(n89),
	.A2(write),
	.A1(data[12]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U28 (
	.ZN(n56),
	.B2(n72),
	.B1(FE_OFN28_write),
	.A(n88), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U29 (
	.ZN(n88),
	.A2(FE_OFN28_write),
	.A1(data[13]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U30 (
	.ZN(n55),
	.B2(n71),
	.B1(write),
	.A(n87), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U31 (
	.ZN(n87),
	.A2(write),
	.A1(data[14]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U32 (
	.ZN(n54),
	.A(reset), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U33 (
	.ZN(n53),
	.B2(n70),
	.B1(write),
	.A(n86), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U34 (
	.ZN(n86),
	.A2(write),
	.A1(data[15]), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module SingleReg_12 (
	data, 
	clk, 
	reset, 
	write, 
	dataOut, 
	FE_OFN12_write, 
	FE_OFN3_write, 
	FE_OFN23_write, 
	FE_OFN26_write, 
	FE_OFN28_write, 
	clk__L2_N8, 
	VDD, 
	VSS);
   input [15:0] data;
   input clk;
   input reset;
   input write;
   output [15:0] dataOut;
   input FE_OFN12_write;
   input FE_OFN3_write;
   input FE_OFN23_write;
   input FE_OFN26_write;
   input FE_OFN28_write;
   input clk__L2_N8;
   inout VDD;
   inout VSS;

   // Internal wires
   wire FE_OFN27_write;
   wire n53;
   wire n54;
   wire n55;
   wire n56;
   wire n57;
   wire n58;
   wire n59;
   wire n60;
   wire n61;
   wire n62;
   wire n63;
   wire n64;
   wire n65;
   wire n66;
   wire n67;
   wire n68;
   wire n69;
   wire n70;
   wire n71;
   wire n72;
   wire n73;
   wire n74;
   wire n75;
   wire n76;
   wire n77;
   wire n78;
   wire n79;
   wire n80;
   wire n81;
   wire n82;
   wire n83;
   wire n84;
   wire n85;
   wire n86;
   wire n87;
   wire n88;
   wire n89;
   wire n90;
   wire n91;
   wire n92;
   wire n93;
   wire n94;
   wire n95;
   wire n96;
   wire n97;
   wire n98;
   wire n99;
   wire n100;
   wire n101;

   // Module instantiations
   BUF_X1 FE_OFC27_write (
	.Z(FE_OFN27_write),
	.A(FE_OFN26_write), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[15]  (
	.RN(n54),
	.QN(n70),
	.Q(dataOut[15]),
	.D(n53),
	.CK(clk__L2_N8), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[14]  (
	.RN(n54),
	.QN(n71),
	.Q(dataOut[14]),
	.D(n55),
	.CK(clk__L2_N8), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[13]  (
	.RN(n54),
	.QN(n72),
	.Q(dataOut[13]),
	.D(n56),
	.CK(clk__L2_N8), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[12]  (
	.RN(n54),
	.QN(n73),
	.Q(dataOut[12]),
	.D(n57),
	.CK(clk__L2_N8), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[11]  (
	.RN(n54),
	.QN(n74),
	.Q(dataOut[11]),
	.D(n58),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[10]  (
	.RN(n54),
	.QN(n75),
	.Q(dataOut[10]),
	.D(n59),
	.CK(clk__L2_N8), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[9]  (
	.RN(n54),
	.QN(n76),
	.Q(dataOut[9]),
	.D(n60),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[8]  (
	.RN(n54),
	.QN(n77),
	.Q(dataOut[8]),
	.D(n61),
	.CK(clk__L2_N8), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[7]  (
	.RN(n54),
	.QN(n78),
	.Q(dataOut[7]),
	.D(n62),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[6]  (
	.RN(n54),
	.QN(n79),
	.Q(dataOut[6]),
	.D(n63),
	.CK(clk__L2_N8), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[5]  (
	.RN(n54),
	.QN(n80),
	.Q(dataOut[5]),
	.D(n64),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[4]  (
	.RN(n54),
	.QN(n81),
	.Q(dataOut[4]),
	.D(n65),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[3]  (
	.RN(n54),
	.QN(n82),
	.Q(dataOut[3]),
	.D(n66),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[2]  (
	.RN(n54),
	.QN(n83),
	.Q(dataOut[2]),
	.D(n67),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[1]  (
	.RN(n54),
	.QN(n84),
	.Q(dataOut[1]),
	.D(n68),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[0]  (
	.RN(n54),
	.QN(n85),
	.Q(dataOut[0]),
	.D(n69),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U2 (
	.ZN(n69),
	.B2(n85),
	.B1(FE_OFN28_write),
	.A(n101), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U3 (
	.ZN(n101),
	.A2(data[0]),
	.A1(FE_OFN28_write), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U4 (
	.ZN(n68),
	.B2(n84),
	.B1(FE_OFN12_write),
	.A(n100), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U5 (
	.ZN(n100),
	.A2(FE_OFN12_write),
	.A1(data[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U6 (
	.ZN(n67),
	.B2(n83),
	.B1(FE_OFN28_write),
	.A(n99), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U7 (
	.ZN(n99),
	.A2(FE_OFN28_write),
	.A1(data[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U8 (
	.ZN(n66),
	.B2(n82),
	.B1(FE_OFN28_write),
	.A(n98), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U9 (
	.ZN(n98),
	.A2(FE_OFN28_write),
	.A1(data[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U10 (
	.ZN(n65),
	.B2(n81),
	.B1(FE_OFN28_write),
	.A(n97), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U11 (
	.ZN(n97),
	.A2(FE_OFN26_write),
	.A1(data[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U12 (
	.ZN(n64),
	.B2(n80),
	.B1(FE_OFN27_write),
	.A(n96), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U13 (
	.ZN(n96),
	.A2(FE_OFN27_write),
	.A1(data[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U14 (
	.ZN(n63),
	.B2(n79),
	.B1(FE_OFN27_write),
	.A(n95), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U15 (
	.ZN(n95),
	.A2(FE_OFN27_write),
	.A1(data[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U16 (
	.ZN(n62),
	.B2(n78),
	.B1(FE_OFN28_write),
	.A(n94), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U17 (
	.ZN(n94),
	.A2(FE_OFN28_write),
	.A1(data[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U18 (
	.ZN(n61),
	.B2(n77),
	.B1(FE_OFN3_write),
	.A(n93), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U19 (
	.ZN(n93),
	.A2(FE_OFN3_write),
	.A1(data[8]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U20 (
	.ZN(n60),
	.B2(n76),
	.B1(FE_OFN28_write),
	.A(n92), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U21 (
	.ZN(n92),
	.A2(FE_OFN26_write),
	.A1(data[9]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U22 (
	.ZN(n59),
	.B2(n75),
	.B1(write),
	.A(n91), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U23 (
	.ZN(n91),
	.A2(write),
	.A1(data[10]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U24 (
	.ZN(n58),
	.B2(n74),
	.B1(FE_OFN3_write),
	.A(n90), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U25 (
	.ZN(n90),
	.A2(FE_OFN3_write),
	.A1(data[11]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U26 (
	.ZN(n57),
	.B2(n73),
	.B1(FE_OFN3_write),
	.A(n89), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U27 (
	.ZN(n89),
	.A2(FE_OFN3_write),
	.A1(data[12]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U28 (
	.ZN(n56),
	.B2(n72),
	.B1(FE_OFN23_write),
	.A(n88), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U29 (
	.ZN(n88),
	.A2(write),
	.A1(data[13]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U30 (
	.ZN(n55),
	.B2(n71),
	.B1(write),
	.A(n87), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U31 (
	.ZN(n87),
	.A2(write),
	.A1(data[14]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U32 (
	.ZN(n54),
	.A(reset), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U33 (
	.ZN(n53),
	.B2(n70),
	.B1(write),
	.A(n86), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U34 (
	.ZN(n86),
	.A2(write),
	.A1(data[15]), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module SingleReg_11 (
	data, 
	clk, 
	reset, 
	write, 
	dataOut, 
	FE_OFN11_write, 
	FE_OFN5_write, 
	FE_OFN8_write, 
	FE_OFN49_write, 
	FE_OFN51_write, 
	FE_OFN53_write, 
	FE_OFN54_write, 
	FE_OFN56_write, 
	clk__L2_N10, 
	clk__L2_N5, 
	clk__L2_N6, 
	VDD, 
	VSS);
   input [15:0] data;
   input clk;
   input reset;
   input write;
   output [15:0] dataOut;
   input FE_OFN11_write;
   input FE_OFN5_write;
   input FE_OFN8_write;
   input FE_OFN49_write;
   input FE_OFN51_write;
   input FE_OFN53_write;
   input FE_OFN54_write;
   input FE_OFN56_write;
   input clk__L2_N10;
   input clk__L2_N5;
   input clk__L2_N6;
   inout VDD;
   inout VSS;

   // Internal wires
   wire n53;
   wire n54;
   wire n55;
   wire n56;
   wire n57;
   wire n58;
   wire n59;
   wire n60;
   wire n61;
   wire n62;
   wire n63;
   wire n64;
   wire n65;
   wire n66;
   wire n67;
   wire n68;
   wire n69;
   wire n70;
   wire n71;
   wire n72;
   wire n73;
   wire n74;
   wire n75;
   wire n76;
   wire n77;
   wire n78;
   wire n79;
   wire n80;
   wire n81;
   wire n82;
   wire n83;
   wire n84;
   wire n85;
   wire n86;
   wire n87;
   wire n88;
   wire n89;
   wire n90;
   wire n91;
   wire n92;
   wire n93;
   wire n94;
   wire n95;
   wire n96;
   wire n97;
   wire n98;
   wire n99;
   wire n100;
   wire n101;

   // Module instantiations
   DFFR_X1 \Reg_reg[15]  (
	.RN(n54),
	.QN(n70),
	.Q(dataOut[15]),
	.D(n53),
	.CK(clk__L2_N6), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[14]  (
	.RN(n54),
	.QN(n71),
	.Q(dataOut[14]),
	.D(n55),
	.CK(clk__L2_N6), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[13]  (
	.RN(n54),
	.QN(n72),
	.Q(dataOut[13]),
	.D(n56),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[12]  (
	.RN(n54),
	.QN(n73),
	.Q(dataOut[12]),
	.D(n57),
	.CK(clk__L2_N5), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[11]  (
	.RN(n54),
	.QN(n74),
	.Q(dataOut[11]),
	.D(n58),
	.CK(clk__L2_N5), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[10]  (
	.RN(n54),
	.QN(n75),
	.Q(dataOut[10]),
	.D(n59),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[9]  (
	.RN(n54),
	.QN(n76),
	.Q(dataOut[9]),
	.D(n60),
	.CK(clk__L2_N10), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[8]  (
	.RN(n54),
	.QN(n77),
	.Q(dataOut[8]),
	.D(n61),
	.CK(clk__L2_N5), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[7]  (
	.RN(n54),
	.QN(n78),
	.Q(dataOut[7]),
	.D(n62),
	.CK(clk__L2_N5), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[6]  (
	.RN(n54),
	.QN(n79),
	.Q(dataOut[6]),
	.D(n63),
	.CK(clk__L2_N5), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[5]  (
	.RN(n54),
	.QN(n80),
	.Q(dataOut[5]),
	.D(n64),
	.CK(clk__L2_N10), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[4]  (
	.RN(n54),
	.QN(n81),
	.Q(dataOut[4]),
	.D(n65),
	.CK(clk__L2_N5), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[3]  (
	.RN(n54),
	.QN(n82),
	.Q(dataOut[3]),
	.D(n66),
	.CK(clk__L2_N5), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[2]  (
	.RN(n54),
	.QN(n83),
	.Q(dataOut[2]),
	.D(n67),
	.CK(clk__L2_N5), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[1]  (
	.RN(n54),
	.QN(n84),
	.Q(dataOut[1]),
	.D(n68),
	.CK(clk__L2_N5), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[0]  (
	.RN(n54),
	.QN(n85),
	.Q(dataOut[0]),
	.D(n69),
	.CK(clk__L2_N5), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U2 (
	.ZN(n69),
	.B2(n85),
	.B1(write),
	.A(n101), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U3 (
	.ZN(n101),
	.A2(data[0]),
	.A1(write), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U4 (
	.ZN(n68),
	.B2(n84),
	.B1(FE_OFN56_write),
	.A(n100), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U5 (
	.ZN(n100),
	.A2(FE_OFN56_write),
	.A1(data[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U6 (
	.ZN(n67),
	.B2(n83),
	.B1(FE_OFN56_write),
	.A(n99), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U7 (
	.ZN(n99),
	.A2(FE_OFN56_write),
	.A1(data[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U8 (
	.ZN(n66),
	.B2(n82),
	.B1(FE_OFN56_write),
	.A(n98), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U9 (
	.ZN(n98),
	.A2(FE_OFN56_write),
	.A1(data[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U10 (
	.ZN(n65),
	.B2(n81),
	.B1(FE_OFN54_write),
	.A(n97), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U11 (
	.ZN(n97),
	.A2(FE_OFN11_write),
	.A1(data[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U12 (
	.ZN(n64),
	.B2(n80),
	.B1(FE_OFN54_write),
	.A(n96), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U13 (
	.ZN(n96),
	.A2(FE_OFN54_write),
	.A1(data[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U14 (
	.ZN(n63),
	.B2(n79),
	.B1(FE_OFN11_write),
	.A(n95), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U15 (
	.ZN(n95),
	.A2(FE_OFN11_write),
	.A1(data[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U16 (
	.ZN(n62),
	.B2(n78),
	.B1(write),
	.A(n94), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U17 (
	.ZN(n94),
	.A2(write),
	.A1(data[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U18 (
	.ZN(n61),
	.B2(n77),
	.B1(FE_OFN49_write),
	.A(n93), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U19 (
	.ZN(n93),
	.A2(FE_OFN49_write),
	.A1(data[8]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U20 (
	.ZN(n60),
	.B2(n76),
	.B1(write),
	.A(n92), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U21 (
	.ZN(n92),
	.A2(write),
	.A1(data[9]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U22 (
	.ZN(n59),
	.B2(n75),
	.B1(FE_OFN49_write),
	.A(n91), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U23 (
	.ZN(n91),
	.A2(FE_OFN8_write),
	.A1(data[10]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U24 (
	.ZN(n58),
	.B2(n74),
	.B1(FE_OFN11_write),
	.A(n90), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U25 (
	.ZN(n90),
	.A2(FE_OFN11_write),
	.A1(data[11]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U26 (
	.ZN(n57),
	.B2(n73),
	.B1(FE_OFN5_write),
	.A(n89), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U27 (
	.ZN(n89),
	.A2(FE_OFN53_write),
	.A1(data[12]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U28 (
	.ZN(n56),
	.B2(n72),
	.B1(FE_OFN49_write),
	.A(n88), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U29 (
	.ZN(n88),
	.A2(FE_OFN49_write),
	.A1(data[13]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U30 (
	.ZN(n55),
	.B2(n71),
	.B1(FE_OFN5_write),
	.A(n87), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U31 (
	.ZN(n87),
	.A2(FE_OFN5_write),
	.A1(data[14]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X2 U32 (
	.ZN(n54),
	.A(reset), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U33 (
	.ZN(n53),
	.B2(n70),
	.B1(FE_OFN51_write),
	.A(n86), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U34 (
	.ZN(n86),
	.A2(FE_OFN51_write),
	.A1(data[15]), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module SingleReg_10 (
	data, 
	clk, 
	reset, 
	write, 
	dataOut, 
	FE_OFN11_write, 
	FE_OFN4_write, 
	FE_OFN5_write, 
	FE_OFN8_write, 
	FE_OFN48_write, 
	FE_OFN49_write, 
	FE_OFN54_write, 
	FE_OFN56_write, 
	clk__L2_N10, 
	clk__L2_N5, 
	VDD, 
	VSS);
   input [15:0] data;
   input clk;
   input reset;
   input write;
   output [15:0] dataOut;
   input FE_OFN11_write;
   input FE_OFN4_write;
   input FE_OFN5_write;
   input FE_OFN8_write;
   input FE_OFN48_write;
   input FE_OFN49_write;
   input FE_OFN54_write;
   input FE_OFN56_write;
   input clk__L2_N10;
   input clk__L2_N5;
   inout VDD;
   inout VSS;

   // Internal wires
   wire n53;
   wire n54;
   wire n55;
   wire n56;
   wire n57;
   wire n58;
   wire n59;
   wire n60;
   wire n61;
   wire n62;
   wire n63;
   wire n64;
   wire n65;
   wire n66;
   wire n67;
   wire n68;
   wire n69;
   wire n70;
   wire n71;
   wire n72;
   wire n73;
   wire n74;
   wire n75;
   wire n76;
   wire n77;
   wire n78;
   wire n79;
   wire n80;
   wire n81;
   wire n82;
   wire n83;
   wire n84;
   wire n85;
   wire n86;
   wire n87;
   wire n88;
   wire n89;
   wire n90;
   wire n91;
   wire n92;
   wire n93;
   wire n94;
   wire n95;
   wire n96;
   wire n97;
   wire n98;
   wire n99;
   wire n100;
   wire n101;

   // Module instantiations
   DFFR_X1 \Reg_reg[15]  (
	.RN(n54),
	.QN(n70),
	.Q(dataOut[15]),
	.D(n53),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[14]  (
	.RN(n54),
	.QN(n71),
	.Q(dataOut[14]),
	.D(n55),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[13]  (
	.RN(n54),
	.QN(n72),
	.Q(dataOut[13]),
	.D(n56),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[12]  (
	.RN(n54),
	.QN(n73),
	.Q(dataOut[12]),
	.D(n57),
	.CK(clk__L2_N5), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[11]  (
	.RN(n54),
	.QN(n74),
	.Q(dataOut[11]),
	.D(n58),
	.CK(clk__L2_N5), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[10]  (
	.RN(n54),
	.QN(n75),
	.Q(dataOut[10]),
	.D(n59),
	.CK(clk__L2_N5), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[9]  (
	.RN(n54),
	.QN(n76),
	.Q(dataOut[9]),
	.D(n60),
	.CK(clk__L2_N10), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[8]  (
	.RN(n54),
	.QN(n77),
	.Q(dataOut[8]),
	.D(n61),
	.CK(clk__L2_N5), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[7]  (
	.RN(n54),
	.QN(n78),
	.Q(dataOut[7]),
	.D(n62),
	.CK(clk__L2_N10), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[6]  (
	.RN(n54),
	.QN(n79),
	.Q(dataOut[6]),
	.D(n63),
	.CK(clk__L2_N5), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[5]  (
	.RN(n54),
	.QN(n80),
	.Q(dataOut[5]),
	.D(n64),
	.CK(clk__L2_N5), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[4]  (
	.RN(n54),
	.QN(n81),
	.Q(dataOut[4]),
	.D(n65),
	.CK(clk__L2_N5), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[3]  (
	.RN(n54),
	.QN(n82),
	.Q(dataOut[3]),
	.D(n66),
	.CK(clk__L2_N5), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[2]  (
	.RN(n54),
	.QN(n83),
	.Q(dataOut[2]),
	.D(n67),
	.CK(clk__L2_N5), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[1]  (
	.RN(n54),
	.QN(n84),
	.Q(dataOut[1]),
	.D(n68),
	.CK(clk__L2_N5), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[0]  (
	.RN(n54),
	.QN(n85),
	.Q(dataOut[0]),
	.D(n69),
	.CK(clk__L2_N5), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U2 (
	.ZN(n69),
	.B2(n85),
	.B1(FE_OFN48_write),
	.A(n101), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U3 (
	.ZN(n101),
	.A2(data[0]),
	.A1(FE_OFN48_write), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U4 (
	.ZN(n68),
	.B2(n84),
	.B1(FE_OFN56_write),
	.A(n100), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U5 (
	.ZN(n100),
	.A2(FE_OFN56_write),
	.A1(data[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U6 (
	.ZN(n67),
	.B2(n83),
	.B1(FE_OFN48_write),
	.A(n99), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U7 (
	.ZN(n99),
	.A2(FE_OFN48_write),
	.A1(data[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U8 (
	.ZN(n66),
	.B2(n82),
	.B1(FE_OFN48_write),
	.A(n98), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U9 (
	.ZN(n98),
	.A2(FE_OFN48_write),
	.A1(data[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U10 (
	.ZN(n65),
	.B2(n81),
	.B1(FE_OFN11_write),
	.A(n97), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U11 (
	.ZN(n97),
	.A2(FE_OFN11_write),
	.A1(data[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U12 (
	.ZN(n64),
	.B2(n80),
	.B1(write),
	.A(n96), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U13 (
	.ZN(n96),
	.A2(FE_OFN54_write),
	.A1(data[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U14 (
	.ZN(n63),
	.B2(n79),
	.B1(FE_OFN54_write),
	.A(n95), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U15 (
	.ZN(n95),
	.A2(FE_OFN11_write),
	.A1(data[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U16 (
	.ZN(n62),
	.B2(n78),
	.B1(FE_OFN48_write),
	.A(n94), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U17 (
	.ZN(n94),
	.A2(FE_OFN48_write),
	.A1(data[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U18 (
	.ZN(n61),
	.B2(n77),
	.B1(FE_OFN8_write),
	.A(n93), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U19 (
	.ZN(n93),
	.A2(FE_OFN8_write),
	.A1(data[8]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U20 (
	.ZN(n60),
	.B2(n76),
	.B1(FE_OFN48_write),
	.A(n92), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U21 (
	.ZN(n92),
	.A2(FE_OFN48_write),
	.A1(data[9]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U22 (
	.ZN(n59),
	.B2(n75),
	.B1(FE_OFN49_write),
	.A(n91), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U23 (
	.ZN(n91),
	.A2(FE_OFN49_write),
	.A1(data[10]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U24 (
	.ZN(n58),
	.B2(n74),
	.B1(FE_OFN11_write),
	.A(n90), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U25 (
	.ZN(n90),
	.A2(FE_OFN11_write),
	.A1(data[11]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U26 (
	.ZN(n57),
	.B2(n73),
	.B1(FE_OFN5_write),
	.A(n89), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U27 (
	.ZN(n89),
	.A2(FE_OFN5_write),
	.A1(data[12]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U28 (
	.ZN(n56),
	.B2(n72),
	.B1(FE_OFN49_write),
	.A(n88), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U29 (
	.ZN(n88),
	.A2(FE_OFN49_write),
	.A1(data[13]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U30 (
	.ZN(n55),
	.B2(n71),
	.B1(FE_OFN4_write),
	.A(n87), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U31 (
	.ZN(n87),
	.A2(FE_OFN4_write),
	.A1(data[14]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X2 U32 (
	.ZN(n54),
	.A(reset), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U33 (
	.ZN(n53),
	.B2(n70),
	.B1(FE_OFN5_write),
	.A(n86), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U34 (
	.ZN(n86),
	.A2(FE_OFN5_write),
	.A1(data[15]), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module SingleReg_9 (
	data, 
	clk, 
	reset, 
	write, 
	dataOut, 
	FE_OFN13_write, 
	FE_OFN5_write, 
	FE_OFN56_write, 
	FE_OFN57_write, 
	FE_OFN58_write, 
	clk__L2_N6, 
	clk__L2_N9, 
	VDD, 
	VSS);
   input [15:0] data;
   input clk;
   input reset;
   input write;
   output [15:0] dataOut;
   input FE_OFN13_write;
   input FE_OFN5_write;
   input FE_OFN56_write;
   input FE_OFN57_write;
   input FE_OFN58_write;
   input clk__L2_N6;
   input clk__L2_N9;
   inout VDD;
   inout VSS;

   // Internal wires
   wire n53;
   wire n54;
   wire n55;
   wire n56;
   wire n57;
   wire n58;
   wire n59;
   wire n60;
   wire n61;
   wire n62;
   wire n63;
   wire n64;
   wire n65;
   wire n66;
   wire n67;
   wire n68;
   wire n69;
   wire n70;
   wire n71;
   wire n72;
   wire n73;
   wire n74;
   wire n75;
   wire n76;
   wire n77;
   wire n78;
   wire n79;
   wire n80;
   wire n81;
   wire n82;
   wire n83;
   wire n84;
   wire n85;
   wire n86;
   wire n87;
   wire n88;
   wire n89;
   wire n90;
   wire n91;
   wire n92;
   wire n93;
   wire n94;
   wire n95;
   wire n96;
   wire n97;
   wire n98;
   wire n99;
   wire n100;
   wire n101;

   // Module instantiations
   DFFR_X1 \Reg_reg[15]  (
	.RN(n54),
	.QN(n70),
	.Q(dataOut[15]),
	.D(n53),
	.CK(clk__L2_N6), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[14]  (
	.RN(n54),
	.QN(n71),
	.Q(dataOut[14]),
	.D(n55),
	.CK(clk__L2_N6), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[13]  (
	.RN(n54),
	.QN(n72),
	.Q(dataOut[13]),
	.D(n56),
	.CK(clk__L2_N6), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[12]  (
	.RN(n54),
	.QN(n73),
	.Q(dataOut[12]),
	.D(n57),
	.CK(clk__L2_N6), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[11]  (
	.RN(n54),
	.QN(n74),
	.Q(dataOut[11]),
	.D(n58),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[10]  (
	.RN(n54),
	.QN(n75),
	.Q(dataOut[10]),
	.D(n59),
	.CK(clk__L2_N6), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[9]  (
	.RN(n54),
	.QN(n76),
	.Q(dataOut[9]),
	.D(n60),
	.CK(clk__L2_N9), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[8]  (
	.RN(n54),
	.QN(n77),
	.Q(dataOut[8]),
	.D(n61),
	.CK(clk__L2_N6), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[7]  (
	.RN(n54),
	.QN(n78),
	.Q(dataOut[7]),
	.D(n62),
	.CK(clk__L2_N9), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[6]  (
	.RN(n54),
	.QN(n79),
	.Q(dataOut[6]),
	.D(n63),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[5]  (
	.RN(n54),
	.QN(n80),
	.Q(dataOut[5]),
	.D(n64),
	.CK(clk__L2_N9), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[4]  (
	.RN(n54),
	.QN(n81),
	.Q(dataOut[4]),
	.D(n65),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[3]  (
	.RN(n54),
	.QN(n82),
	.Q(dataOut[3]),
	.D(n66),
	.CK(clk__L2_N9), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[2]  (
	.RN(n54),
	.QN(n83),
	.Q(dataOut[2]),
	.D(n67),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[1]  (
	.RN(n54),
	.QN(n84),
	.Q(dataOut[1]),
	.D(n68),
	.CK(clk__L2_N9), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[0]  (
	.RN(n54),
	.QN(n85),
	.Q(dataOut[0]),
	.D(n69),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U2 (
	.ZN(n69),
	.B2(n85),
	.B1(FE_OFN56_write),
	.A(n101), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U3 (
	.ZN(n101),
	.A2(data[0]),
	.A1(FE_OFN56_write), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U4 (
	.ZN(n68),
	.B2(n84),
	.B1(FE_OFN56_write),
	.A(n100), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U5 (
	.ZN(n100),
	.A2(FE_OFN56_write),
	.A1(data[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U6 (
	.ZN(n67),
	.B2(n83),
	.B1(FE_OFN56_write),
	.A(n99), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U7 (
	.ZN(n99),
	.A2(FE_OFN56_write),
	.A1(data[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U8 (
	.ZN(n66),
	.B2(n82),
	.B1(FE_OFN56_write),
	.A(n98), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U9 (
	.ZN(n98),
	.A2(FE_OFN56_write),
	.A1(data[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U10 (
	.ZN(n65),
	.B2(n81),
	.B1(write),
	.A(n97), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U11 (
	.ZN(n97),
	.A2(write),
	.A1(data[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U12 (
	.ZN(n64),
	.B2(n80),
	.B1(FE_OFN13_write),
	.A(n96), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U13 (
	.ZN(n96),
	.A2(FE_OFN57_write),
	.A1(data[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U14 (
	.ZN(n63),
	.B2(n79),
	.B1(FE_OFN13_write),
	.A(n95), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U15 (
	.ZN(n95),
	.A2(FE_OFN13_write),
	.A1(data[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U16 (
	.ZN(n62),
	.B2(n78),
	.B1(FE_OFN56_write),
	.A(n94), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U17 (
	.ZN(n94),
	.A2(FE_OFN56_write),
	.A1(data[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U18 (
	.ZN(n61),
	.B2(n77),
	.B1(FE_OFN57_write),
	.A(n93), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U19 (
	.ZN(n93),
	.A2(FE_OFN57_write),
	.A1(data[8]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U20 (
	.ZN(n60),
	.B2(n76),
	.B1(FE_OFN58_write),
	.A(n92), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U21 (
	.ZN(n92),
	.A2(FE_OFN58_write),
	.A1(data[9]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U22 (
	.ZN(n59),
	.B2(n75),
	.B1(FE_OFN57_write),
	.A(n91), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U23 (
	.ZN(n91),
	.A2(FE_OFN57_write),
	.A1(data[10]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U24 (
	.ZN(n58),
	.B2(n74),
	.B1(FE_OFN57_write),
	.A(n90), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U25 (
	.ZN(n90),
	.A2(FE_OFN57_write),
	.A1(data[11]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U26 (
	.ZN(n57),
	.B2(n73),
	.B1(FE_OFN5_write),
	.A(n89), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U27 (
	.ZN(n89),
	.A2(FE_OFN5_write),
	.A1(data[12]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U28 (
	.ZN(n56),
	.B2(n72),
	.B1(FE_OFN57_write),
	.A(n88), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U29 (
	.ZN(n88),
	.A2(FE_OFN5_write),
	.A1(data[13]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U30 (
	.ZN(n55),
	.B2(n71),
	.B1(FE_OFN5_write),
	.A(n87), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U31 (
	.ZN(n87),
	.A2(FE_OFN5_write),
	.A1(data[14]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U32 (
	.ZN(n54),
	.A(reset), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U33 (
	.ZN(n53),
	.B2(n70),
	.B1(FE_OFN5_write),
	.A(n86), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U34 (
	.ZN(n86),
	.A2(FE_OFN5_write),
	.A1(data[15]), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module SingleReg_8 (
	data, 
	clk, 
	reset, 
	write, 
	dataOut, 
	FE_OFN13_write, 
	FE_OFN5_write, 
	FE_OFN8_write, 
	FE_OFN53_write, 
	FE_OFN54_write, 
	FE_OFN56_write, 
	clk__L2_N5, 
	clk__L2_N6, 
	VDD, 
	VSS);
   input [15:0] data;
   input clk;
   input reset;
   input write;
   output [15:0] dataOut;
   input FE_OFN13_write;
   input FE_OFN5_write;
   input FE_OFN8_write;
   input FE_OFN53_write;
   input FE_OFN54_write;
   input FE_OFN56_write;
   input clk__L2_N5;
   input clk__L2_N6;
   inout VDD;
   inout VSS;

   // Internal wires
   wire n53;
   wire n54;
   wire n55;
   wire n56;
   wire n57;
   wire n58;
   wire n59;
   wire n60;
   wire n61;
   wire n62;
   wire n63;
   wire n64;
   wire n65;
   wire n66;
   wire n67;
   wire n68;
   wire n69;
   wire n70;
   wire n71;
   wire n72;
   wire n73;
   wire n74;
   wire n75;
   wire n76;
   wire n77;
   wire n78;
   wire n79;
   wire n80;
   wire n81;
   wire n82;
   wire n83;
   wire n84;
   wire n85;
   wire n86;
   wire n87;
   wire n88;
   wire n89;
   wire n90;
   wire n91;
   wire n92;
   wire n93;
   wire n94;
   wire n95;
   wire n96;
   wire n97;
   wire n98;
   wire n99;
   wire n100;
   wire n101;

   // Module instantiations
   DFFR_X1 \Reg_reg[15]  (
	.RN(n54),
	.QN(n70),
	.Q(dataOut[15]),
	.D(n53),
	.CK(clk__L2_N6), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[14]  (
	.RN(n54),
	.QN(n71),
	.Q(dataOut[14]),
	.D(n55),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[13]  (
	.RN(n54),
	.QN(n72),
	.Q(dataOut[13]),
	.D(n56),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[12]  (
	.RN(n54),
	.QN(n73),
	.Q(dataOut[12]),
	.D(n57),
	.CK(clk__L2_N5), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[11]  (
	.RN(n54),
	.QN(n74),
	.Q(dataOut[11]),
	.D(n58),
	.CK(clk__L2_N5), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[10]  (
	.RN(n54),
	.QN(n75),
	.Q(dataOut[10]),
	.D(n59),
	.CK(clk__L2_N6), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[9]  (
	.RN(n54),
	.QN(n76),
	.Q(dataOut[9]),
	.D(n60),
	.CK(clk__L2_N5), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[8]  (
	.RN(n54),
	.QN(n77),
	.Q(dataOut[8]),
	.D(n61),
	.CK(clk__L2_N6), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[7]  (
	.RN(n54),
	.QN(n78),
	.Q(dataOut[7]),
	.D(n62),
	.CK(clk__L2_N5), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[6]  (
	.RN(n54),
	.QN(n79),
	.Q(dataOut[6]),
	.D(n63),
	.CK(clk__L2_N5), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[5]  (
	.RN(n54),
	.QN(n80),
	.Q(dataOut[5]),
	.D(n64),
	.CK(clk__L2_N5), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[4]  (
	.RN(n54),
	.QN(n81),
	.Q(dataOut[4]),
	.D(n65),
	.CK(clk__L2_N5), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[3]  (
	.RN(n54),
	.QN(n82),
	.Q(dataOut[3]),
	.D(n66),
	.CK(clk__L2_N5), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[2]  (
	.RN(n54),
	.QN(n83),
	.Q(dataOut[2]),
	.D(n67),
	.CK(clk__L2_N5), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[1]  (
	.RN(n54),
	.QN(n84),
	.Q(dataOut[1]),
	.D(n68),
	.CK(clk__L2_N5), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[0]  (
	.RN(n54),
	.QN(n85),
	.Q(dataOut[0]),
	.D(n69),
	.CK(clk__L2_N5), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U2 (
	.ZN(n69),
	.B2(n85),
	.B1(write),
	.A(n101), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U3 (
	.ZN(n101),
	.A2(data[0]),
	.A1(write), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U4 (
	.ZN(n68),
	.B2(n84),
	.B1(FE_OFN56_write),
	.A(n100), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U5 (
	.ZN(n100),
	.A2(FE_OFN56_write),
	.A1(data[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U6 (
	.ZN(n67),
	.B2(n83),
	.B1(FE_OFN56_write),
	.A(n99), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U7 (
	.ZN(n99),
	.A2(FE_OFN56_write),
	.A1(data[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U8 (
	.ZN(n66),
	.B2(n82),
	.B1(FE_OFN56_write),
	.A(n98), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U9 (
	.ZN(n98),
	.A2(write),
	.A1(data[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U10 (
	.ZN(n65),
	.B2(n81),
	.B1(write),
	.A(n97), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U11 (
	.ZN(n97),
	.A2(write),
	.A1(data[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U12 (
	.ZN(n64),
	.B2(n80),
	.B1(FE_OFN8_write),
	.A(n96), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U13 (
	.ZN(n96),
	.A2(FE_OFN8_write),
	.A1(data[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U14 (
	.ZN(n63),
	.B2(n79),
	.B1(write),
	.A(n95), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U15 (
	.ZN(n95),
	.A2(FE_OFN13_write),
	.A1(data[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U16 (
	.ZN(n62),
	.B2(n78),
	.B1(write),
	.A(n94), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U17 (
	.ZN(n94),
	.A2(write),
	.A1(data[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U18 (
	.ZN(n61),
	.B2(n77),
	.B1(FE_OFN13_write),
	.A(n93), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U19 (
	.ZN(n93),
	.A2(FE_OFN13_write),
	.A1(data[8]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U20 (
	.ZN(n60),
	.B2(n76),
	.B1(FE_OFN54_write),
	.A(n92), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U21 (
	.ZN(n92),
	.A2(FE_OFN54_write),
	.A1(data[9]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U22 (
	.ZN(n59),
	.B2(n75),
	.B1(FE_OFN53_write),
	.A(n91), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U23 (
	.ZN(n91),
	.A2(FE_OFN53_write),
	.A1(data[10]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U24 (
	.ZN(n58),
	.B2(n74),
	.B1(FE_OFN53_write),
	.A(n90), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U25 (
	.ZN(n90),
	.A2(FE_OFN13_write),
	.A1(data[11]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U26 (
	.ZN(n57),
	.B2(n73),
	.B1(FE_OFN53_write),
	.A(n89), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U27 (
	.ZN(n89),
	.A2(FE_OFN53_write),
	.A1(data[12]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U28 (
	.ZN(n56),
	.B2(n72),
	.B1(FE_OFN5_write),
	.A(n88), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U29 (
	.ZN(n88),
	.A2(FE_OFN5_write),
	.A1(data[13]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U30 (
	.ZN(n55),
	.B2(n71),
	.B1(FE_OFN5_write),
	.A(n87), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U31 (
	.ZN(n87),
	.A2(FE_OFN5_write),
	.A1(data[14]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U32 (
	.ZN(n54),
	.A(reset), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U33 (
	.ZN(n53),
	.B2(n70),
	.B1(FE_OFN5_write),
	.A(n86), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U34 (
	.ZN(n86),
	.A2(FE_OFN5_write),
	.A1(data[15]), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module SingleReg_7 (
	data, 
	clk, 
	reset, 
	write, 
	dataOut, 
	FE_OFN11_write, 
	FE_OFN5_write, 
	FE_OFN8_write, 
	FE_OFN42_write, 
	FE_OFN46_write, 
	FE_OFN48_write, 
	clk__L2_N10, 
	clk__L2_N4, 
	VDD, 
	VSS);
   input [15:0] data;
   input clk;
   input reset;
   input write;
   output [15:0] dataOut;
   input FE_OFN11_write;
   input FE_OFN5_write;
   input FE_OFN8_write;
   input FE_OFN42_write;
   input FE_OFN46_write;
   input FE_OFN48_write;
   input clk__L2_N10;
   input clk__L2_N4;
   inout VDD;
   inout VSS;

   // Internal wires
   wire n53;
   wire n54;
   wire n55;
   wire n56;
   wire n57;
   wire n58;
   wire n59;
   wire n60;
   wire n61;
   wire n62;
   wire n63;
   wire n64;
   wire n65;
   wire n66;
   wire n67;
   wire n68;
   wire n69;
   wire n70;
   wire n71;
   wire n72;
   wire n73;
   wire n74;
   wire n75;
   wire n76;
   wire n77;
   wire n78;
   wire n79;
   wire n80;
   wire n81;
   wire n82;
   wire n83;
   wire n84;
   wire n85;
   wire n86;
   wire n87;
   wire n88;
   wire n89;
   wire n90;
   wire n91;
   wire n92;
   wire n93;
   wire n94;
   wire n95;
   wire n96;
   wire n97;
   wire n98;
   wire n99;
   wire n100;
   wire n101;

   // Module instantiations
   DFFR_X1 \Reg_reg[15]  (
	.RN(n54),
	.QN(n70),
	.Q(dataOut[15]),
	.D(n53),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[14]  (
	.RN(n54),
	.QN(n71),
	.Q(dataOut[14]),
	.D(n55),
	.CK(clk__L2_N4), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[13]  (
	.RN(n54),
	.QN(n72),
	.Q(dataOut[13]),
	.D(n56),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[12]  (
	.RN(n54),
	.QN(n73),
	.Q(dataOut[12]),
	.D(n57),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[11]  (
	.RN(n54),
	.QN(n74),
	.Q(dataOut[11]),
	.D(n58),
	.CK(clk__L2_N4), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[10]  (
	.RN(n54),
	.QN(n75),
	.Q(dataOut[10]),
	.D(n59),
	.CK(clk__L2_N4), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[9]  (
	.RN(n54),
	.QN(n76),
	.Q(dataOut[9]),
	.D(n60),
	.CK(clk__L2_N10), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[8]  (
	.RN(n54),
	.QN(n77),
	.Q(dataOut[8]),
	.D(n61),
	.CK(clk__L2_N10), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[7]  (
	.RN(n54),
	.QN(n78),
	.Q(dataOut[7]),
	.D(n62),
	.CK(clk__L2_N10), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[6]  (
	.RN(n54),
	.QN(n79),
	.Q(dataOut[6]),
	.D(n63),
	.CK(clk__L2_N10), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[5]  (
	.RN(n54),
	.QN(n80),
	.Q(dataOut[5]),
	.D(n64),
	.CK(clk__L2_N10), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[4]  (
	.RN(n54),
	.QN(n81),
	.Q(dataOut[4]),
	.D(n65),
	.CK(clk__L2_N10), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[3]  (
	.RN(n54),
	.QN(n82),
	.Q(dataOut[3]),
	.D(n66),
	.CK(clk__L2_N10), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[2]  (
	.RN(n54),
	.QN(n83),
	.Q(dataOut[2]),
	.D(n67),
	.CK(clk__L2_N10), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[1]  (
	.RN(n54),
	.QN(n84),
	.Q(dataOut[1]),
	.D(n68),
	.CK(clk__L2_N10), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[0]  (
	.RN(n54),
	.QN(n85),
	.Q(dataOut[0]),
	.D(n69),
	.CK(clk__L2_N10), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U2 (
	.ZN(n69),
	.B2(n85),
	.B1(FE_OFN46_write),
	.A(n101), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U3 (
	.ZN(n101),
	.A2(data[0]),
	.A1(FE_OFN46_write), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U4 (
	.ZN(n68),
	.B2(n84),
	.B1(write),
	.A(n100), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U5 (
	.ZN(n100),
	.A2(write),
	.A1(data[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U6 (
	.ZN(n67),
	.B2(n83),
	.B1(FE_OFN48_write),
	.A(n99), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U7 (
	.ZN(n99),
	.A2(FE_OFN46_write),
	.A1(data[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U8 (
	.ZN(n66),
	.B2(n82),
	.B1(FE_OFN46_write),
	.A(n98), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U9 (
	.ZN(n98),
	.A2(FE_OFN46_write),
	.A1(data[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U10 (
	.ZN(n65),
	.B2(n81),
	.B1(FE_OFN11_write),
	.A(n97), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U11 (
	.ZN(n97),
	.A2(FE_OFN11_write),
	.A1(data[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U12 (
	.ZN(n64),
	.B2(n80),
	.B1(FE_OFN46_write),
	.A(n96), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U13 (
	.ZN(n96),
	.A2(FE_OFN46_write),
	.A1(data[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U14 (
	.ZN(n63),
	.B2(n79),
	.B1(FE_OFN42_write),
	.A(n95), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U15 (
	.ZN(n95),
	.A2(FE_OFN42_write),
	.A1(data[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U16 (
	.ZN(n62),
	.B2(n78),
	.B1(FE_OFN11_write),
	.A(n94), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U17 (
	.ZN(n94),
	.A2(write),
	.A1(data[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U18 (
	.ZN(n61),
	.B2(n77),
	.B1(FE_OFN8_write),
	.A(n93), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U19 (
	.ZN(n93),
	.A2(FE_OFN8_write),
	.A1(data[8]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U20 (
	.ZN(n60),
	.B2(n76),
	.B1(FE_OFN46_write),
	.A(n92), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U21 (
	.ZN(n92),
	.A2(FE_OFN46_write),
	.A1(data[9]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U22 (
	.ZN(n59),
	.B2(n75),
	.B1(FE_OFN5_write),
	.A(n91), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U23 (
	.ZN(n91),
	.A2(FE_OFN5_write),
	.A1(data[10]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U24 (
	.ZN(n58),
	.B2(n74),
	.B1(FE_OFN42_write),
	.A(n90), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U25 (
	.ZN(n90),
	.A2(FE_OFN8_write),
	.A1(data[11]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U26 (
	.ZN(n57),
	.B2(n73),
	.B1(FE_OFN5_write),
	.A(n89), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U27 (
	.ZN(n89),
	.A2(FE_OFN5_write),
	.A1(data[12]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U28 (
	.ZN(n56),
	.B2(n72),
	.B1(FE_OFN5_write),
	.A(n88), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U29 (
	.ZN(n88),
	.A2(FE_OFN5_write),
	.A1(data[13]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U30 (
	.ZN(n55),
	.B2(n71),
	.B1(FE_OFN5_write),
	.A(n87), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U31 (
	.ZN(n87),
	.A2(FE_OFN5_write),
	.A1(data[14]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U32 (
	.ZN(n54),
	.A(reset), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U33 (
	.ZN(n53),
	.B2(n70),
	.B1(FE_OFN5_write),
	.A(n86), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U34 (
	.ZN(n86),
	.A2(FE_OFN5_write),
	.A1(data[15]), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module SingleReg_6 (
	data, 
	clk, 
	reset, 
	write, 
	dataOut, 
	FE_OFN5_write, 
	FE_OFN8_write, 
	FE_OFN42_write, 
	FE_OFN46_write, 
	FE_OFN48_write, 
	clk__L2_N10, 
	clk__L2_N4, 
	VDD, 
	VSS);
   input [15:0] data;
   input clk;
   input reset;
   input write;
   output [15:0] dataOut;
   input FE_OFN5_write;
   input FE_OFN8_write;
   input FE_OFN42_write;
   input FE_OFN46_write;
   input FE_OFN48_write;
   input clk__L2_N10;
   input clk__L2_N4;
   inout VDD;
   inout VSS;

   // Internal wires
   wire n53;
   wire n54;
   wire n55;
   wire n56;
   wire n57;
   wire n58;
   wire n59;
   wire n60;
   wire n61;
   wire n62;
   wire n63;
   wire n64;
   wire n65;
   wire n66;
   wire n67;
   wire n68;
   wire n69;
   wire n70;
   wire n71;
   wire n72;
   wire n73;
   wire n74;
   wire n75;
   wire n76;
   wire n77;
   wire n78;
   wire n79;
   wire n80;
   wire n81;
   wire n82;
   wire n83;
   wire n84;
   wire n85;
   wire n86;
   wire n87;
   wire n88;
   wire n89;
   wire n90;
   wire n91;
   wire n92;
   wire n93;
   wire n94;
   wire n95;
   wire n96;
   wire n97;
   wire n98;
   wire n99;
   wire n100;
   wire n101;

   // Module instantiations
   DFFR_X1 \Reg_reg[15]  (
	.RN(n54),
	.QN(n70),
	.Q(dataOut[15]),
	.D(n53),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[14]  (
	.RN(n54),
	.QN(n71),
	.Q(dataOut[14]),
	.D(n55),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[13]  (
	.RN(n54),
	.QN(n72),
	.Q(dataOut[13]),
	.D(n56),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[12]  (
	.RN(n54),
	.QN(n73),
	.Q(dataOut[12]),
	.D(n57),
	.CK(clk__L2_N4), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[11]  (
	.RN(n54),
	.QN(n74),
	.Q(dataOut[11]),
	.D(n58),
	.CK(clk__L2_N4), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[10]  (
	.RN(n54),
	.QN(n75),
	.Q(dataOut[10]),
	.D(n59),
	.CK(clk__L2_N4), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[9]  (
	.RN(n54),
	.QN(n76),
	.Q(dataOut[9]),
	.D(n60),
	.CK(clk__L2_N10), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[8]  (
	.RN(n54),
	.QN(n77),
	.Q(dataOut[8]),
	.D(n61),
	.CK(clk__L2_N4), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[7]  (
	.RN(n54),
	.QN(n78),
	.Q(dataOut[7]),
	.D(n62),
	.CK(clk__L2_N10), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[6]  (
	.RN(n54),
	.QN(n79),
	.Q(dataOut[6]),
	.D(n63),
	.CK(clk__L2_N10), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[5]  (
	.RN(n54),
	.QN(n80),
	.Q(dataOut[5]),
	.D(n64),
	.CK(clk__L2_N10), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[4]  (
	.RN(n54),
	.QN(n81),
	.Q(dataOut[4]),
	.D(n65),
	.CK(clk__L2_N10), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[3]  (
	.RN(n54),
	.QN(n82),
	.Q(dataOut[3]),
	.D(n66),
	.CK(clk__L2_N10), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[2]  (
	.RN(n54),
	.QN(n83),
	.Q(dataOut[2]),
	.D(n67),
	.CK(clk__L2_N10), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[1]  (
	.RN(n54),
	.QN(n84),
	.Q(dataOut[1]),
	.D(n68),
	.CK(clk__L2_N10), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[0]  (
	.RN(n54),
	.QN(n85),
	.Q(dataOut[0]),
	.D(n69),
	.CK(clk__L2_N10), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U2 (
	.ZN(n69),
	.B2(n85),
	.B1(FE_OFN46_write),
	.A(n101), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U3 (
	.ZN(n101),
	.A2(data[0]),
	.A1(FE_OFN46_write), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U4 (
	.ZN(n68),
	.B2(n84),
	.B1(FE_OFN48_write),
	.A(n100), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U5 (
	.ZN(n100),
	.A2(FE_OFN46_write),
	.A1(data[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U6 (
	.ZN(n67),
	.B2(n83),
	.B1(FE_OFN46_write),
	.A(n99), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U7 (
	.ZN(n99),
	.A2(FE_OFN46_write),
	.A1(data[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U8 (
	.ZN(n66),
	.B2(n82),
	.B1(FE_OFN46_write),
	.A(n98), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U9 (
	.ZN(n98),
	.A2(FE_OFN46_write),
	.A1(data[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U10 (
	.ZN(n65),
	.B2(n81),
	.B1(write),
	.A(n97), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U11 (
	.ZN(n97),
	.A2(write),
	.A1(data[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U12 (
	.ZN(n64),
	.B2(n80),
	.B1(FE_OFN8_write),
	.A(n96), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U13 (
	.ZN(n96),
	.A2(FE_OFN8_write),
	.A1(data[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U14 (
	.ZN(n63),
	.B2(n79),
	.B1(write),
	.A(n95), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U15 (
	.ZN(n95),
	.A2(FE_OFN8_write),
	.A1(data[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U16 (
	.ZN(n62),
	.B2(n78),
	.B1(FE_OFN46_write),
	.A(n94), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U17 (
	.ZN(n94),
	.A2(FE_OFN46_write),
	.A1(data[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U18 (
	.ZN(n61),
	.B2(n77),
	.B1(FE_OFN8_write),
	.A(n93), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U19 (
	.ZN(n93),
	.A2(FE_OFN8_write),
	.A1(data[8]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U20 (
	.ZN(n60),
	.B2(n76),
	.B1(FE_OFN46_write),
	.A(n92), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U21 (
	.ZN(n92),
	.A2(FE_OFN46_write),
	.A1(data[9]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U22 (
	.ZN(n59),
	.B2(n75),
	.B1(FE_OFN8_write),
	.A(n91), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U23 (
	.ZN(n91),
	.A2(FE_OFN8_write),
	.A1(data[10]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U24 (
	.ZN(n58),
	.B2(n74),
	.B1(FE_OFN8_write),
	.A(n90), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U25 (
	.ZN(n90),
	.A2(FE_OFN42_write),
	.A1(data[11]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U26 (
	.ZN(n57),
	.B2(n73),
	.B1(FE_OFN5_write),
	.A(n89), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U27 (
	.ZN(n89),
	.A2(FE_OFN5_write),
	.A1(data[12]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U28 (
	.ZN(n56),
	.B2(n72),
	.B1(FE_OFN5_write),
	.A(n88), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U29 (
	.ZN(n88),
	.A2(FE_OFN5_write),
	.A1(data[13]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U30 (
	.ZN(n55),
	.B2(n71),
	.B1(FE_OFN5_write),
	.A(n87), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U31 (
	.ZN(n87),
	.A2(FE_OFN5_write),
	.A1(data[14]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X2 U32 (
	.ZN(n54),
	.A(reset), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U33 (
	.ZN(n53),
	.B2(n70),
	.B1(FE_OFN5_write),
	.A(n86), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U34 (
	.ZN(n86),
	.A2(FE_OFN5_write),
	.A1(data[15]), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module SingleReg_5 (
	data, 
	clk, 
	reset, 
	write, 
	dataOut, 
	FE_OFN1_write, 
	FE_OFN8_write, 
	FE_OFN35_write, 
	FE_OFN39_write, 
	clk__L2_N4, 
	VDD, 
	VSS);
   input [15:0] data;
   input clk;
   input reset;
   input write;
   output [15:0] dataOut;
   input FE_OFN1_write;
   input FE_OFN8_write;
   input FE_OFN35_write;
   input FE_OFN39_write;
   input clk__L2_N4;
   inout VDD;
   inout VSS;

   // Internal wires
   wire n53;
   wire n54;
   wire n55;
   wire n56;
   wire n57;
   wire n58;
   wire n59;
   wire n60;
   wire n61;
   wire n62;
   wire n63;
   wire n64;
   wire n65;
   wire n66;
   wire n67;
   wire n68;
   wire n69;
   wire n70;
   wire n71;
   wire n72;
   wire n73;
   wire n74;
   wire n75;
   wire n76;
   wire n77;
   wire n78;
   wire n79;
   wire n80;
   wire n81;
   wire n82;
   wire n83;
   wire n84;
   wire n85;
   wire n86;
   wire n87;
   wire n88;
   wire n89;
   wire n90;
   wire n91;
   wire n92;
   wire n93;
   wire n94;
   wire n95;
   wire n96;
   wire n97;
   wire n98;
   wire n99;
   wire n100;
   wire n101;

   // Module instantiations
   DFFR_X1 \Reg_reg[15]  (
	.RN(n54),
	.QN(n70),
	.Q(dataOut[15]),
	.D(n53),
	.CK(clk__L2_N4), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[14]  (
	.RN(n54),
	.QN(n71),
	.Q(dataOut[14]),
	.D(n55),
	.CK(clk__L2_N4), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[13]  (
	.RN(n54),
	.QN(n72),
	.Q(dataOut[13]),
	.D(n56),
	.CK(clk__L2_N4), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[12]  (
	.RN(n54),
	.QN(n73),
	.Q(dataOut[12]),
	.D(n57),
	.CK(clk__L2_N4), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[11]  (
	.RN(n54),
	.QN(n74),
	.Q(dataOut[11]),
	.D(n58),
	.CK(clk__L2_N4), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[10]  (
	.RN(n54),
	.QN(n75),
	.Q(dataOut[10]),
	.D(n59),
	.CK(clk__L2_N4), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[9]  (
	.RN(n54),
	.QN(n76),
	.Q(dataOut[9]),
	.D(n60),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[8]  (
	.RN(n54),
	.QN(n77),
	.Q(dataOut[8]),
	.D(n61),
	.CK(clk__L2_N4), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[7]  (
	.RN(n54),
	.QN(n78),
	.Q(dataOut[7]),
	.D(n62),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[6]  (
	.RN(n54),
	.QN(n79),
	.Q(dataOut[6]),
	.D(n63),
	.CK(clk__L2_N4), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[5]  (
	.RN(n54),
	.QN(n80),
	.Q(dataOut[5]),
	.D(n64),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[4]  (
	.RN(n54),
	.QN(n81),
	.Q(dataOut[4]),
	.D(n65),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[3]  (
	.RN(n54),
	.QN(n82),
	.Q(dataOut[3]),
	.D(n66),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[2]  (
	.RN(n54),
	.QN(n83),
	.Q(dataOut[2]),
	.D(n67),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[1]  (
	.RN(n54),
	.QN(n84),
	.Q(dataOut[1]),
	.D(n68),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[0]  (
	.RN(n54),
	.QN(n85),
	.Q(dataOut[0]),
	.D(n69),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U2 (
	.ZN(n69),
	.B2(n85),
	.B1(write),
	.A(n101), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U3 (
	.ZN(n101),
	.A2(data[0]),
	.A1(write), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U4 (
	.ZN(n68),
	.B2(n84),
	.B1(write),
	.A(n100), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U5 (
	.ZN(n100),
	.A2(write),
	.A1(data[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U6 (
	.ZN(n67),
	.B2(n83),
	.B1(write),
	.A(n99), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U7 (
	.ZN(n99),
	.A2(write),
	.A1(data[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U8 (
	.ZN(n66),
	.B2(n82),
	.B1(write),
	.A(n98), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U9 (
	.ZN(n98),
	.A2(write),
	.A1(data[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U10 (
	.ZN(n65),
	.B2(n81),
	.B1(FE_OFN39_write),
	.A(n97), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U11 (
	.ZN(n97),
	.A2(FE_OFN39_write),
	.A1(data[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U12 (
	.ZN(n64),
	.B2(n80),
	.B1(FE_OFN8_write),
	.A(n96), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U13 (
	.ZN(n96),
	.A2(FE_OFN8_write),
	.A1(data[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U14 (
	.ZN(n63),
	.B2(n79),
	.B1(FE_OFN8_write),
	.A(n95), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U15 (
	.ZN(n95),
	.A2(FE_OFN8_write),
	.A1(data[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U16 (
	.ZN(n62),
	.B2(n78),
	.B1(write),
	.A(n94), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U17 (
	.ZN(n94),
	.A2(write),
	.A1(data[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U18 (
	.ZN(n61),
	.B2(n77),
	.B1(FE_OFN8_write),
	.A(n93), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U19 (
	.ZN(n93),
	.A2(FE_OFN8_write),
	.A1(data[8]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U20 (
	.ZN(n60),
	.B2(n76),
	.B1(write),
	.A(n92), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U21 (
	.ZN(n92),
	.A2(FE_OFN39_write),
	.A1(data[9]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U22 (
	.ZN(n59),
	.B2(n75),
	.B1(FE_OFN8_write),
	.A(n91), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U23 (
	.ZN(n91),
	.A2(FE_OFN8_write),
	.A1(data[10]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U24 (
	.ZN(n58),
	.B2(n74),
	.B1(FE_OFN8_write),
	.A(n90), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U25 (
	.ZN(n90),
	.A2(FE_OFN8_write),
	.A1(data[11]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U26 (
	.ZN(n57),
	.B2(n73),
	.B1(FE_OFN35_write),
	.A(n89), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U27 (
	.ZN(n89),
	.A2(FE_OFN35_write),
	.A1(data[12]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U28 (
	.ZN(n56),
	.B2(n72),
	.B1(FE_OFN35_write),
	.A(n88), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U29 (
	.ZN(n88),
	.A2(FE_OFN35_write),
	.A1(data[13]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U30 (
	.ZN(n55),
	.B2(n71),
	.B1(FE_OFN1_write),
	.A(n87), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U31 (
	.ZN(n87),
	.A2(FE_OFN1_write),
	.A1(data[14]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U32 (
	.ZN(n54),
	.A(reset), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U33 (
	.ZN(n53),
	.B2(n70),
	.B1(FE_OFN1_write),
	.A(n86), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U34 (
	.ZN(n86),
	.A2(FE_OFN35_write),
	.A1(data[15]), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module SingleReg_4 (
	data, 
	clk, 
	reset, 
	write, 
	dataOut, 
	FE_OFN8_write, 
	FE_OFN35_write, 
	FE_OFN39_write, 
	clk__L2_N13, 
	clk__L2_N4, 
	VDD, 
	VSS);
   input [15:0] data;
   input clk;
   input reset;
   input write;
   output [15:0] dataOut;
   input FE_OFN8_write;
   input FE_OFN35_write;
   input FE_OFN39_write;
   input clk__L2_N13;
   input clk__L2_N4;
   inout VDD;
   inout VSS;

   // Internal wires
   wire FE_OFN37_write;
   wire n53;
   wire n54;
   wire n55;
   wire n56;
   wire n57;
   wire n58;
   wire n59;
   wire n60;
   wire n61;
   wire n62;
   wire n63;
   wire n64;
   wire n65;
   wire n66;
   wire n67;
   wire n68;
   wire n69;
   wire n70;
   wire n71;
   wire n72;
   wire n73;
   wire n74;
   wire n75;
   wire n76;
   wire n77;
   wire n78;
   wire n79;
   wire n80;
   wire n81;
   wire n82;
   wire n83;
   wire n84;
   wire n85;
   wire n86;
   wire n87;
   wire n88;
   wire n89;
   wire n90;
   wire n91;
   wire n92;
   wire n93;
   wire n94;
   wire n95;
   wire n96;
   wire n97;
   wire n98;
   wire n99;
   wire n100;
   wire n101;

   // Module instantiations
   BUF_X1 FE_OFC37_write (
	.Z(FE_OFN37_write),
	.A(FE_OFN8_write), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[15]  (
	.RN(n54),
	.QN(n70),
	.Q(dataOut[15]),
	.D(n53),
	.CK(clk__L2_N4), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[14]  (
	.RN(n54),
	.QN(n71),
	.Q(dataOut[14]),
	.D(n55),
	.CK(clk__L2_N4), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[13]  (
	.RN(n54),
	.QN(n72),
	.Q(dataOut[13]),
	.D(n56),
	.CK(clk__L2_N4), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[12]  (
	.RN(n54),
	.QN(n73),
	.Q(dataOut[12]),
	.D(n57),
	.CK(clk__L2_N4), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[11]  (
	.RN(n54),
	.QN(n74),
	.Q(dataOut[11]),
	.D(n58),
	.CK(clk__L2_N4), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[10]  (
	.RN(n54),
	.QN(n75),
	.Q(dataOut[10]),
	.D(n59),
	.CK(clk__L2_N4), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[9]  (
	.RN(n54),
	.QN(n76),
	.Q(dataOut[9]),
	.D(n60),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[8]  (
	.RN(n54),
	.QN(n77),
	.Q(dataOut[8]),
	.D(n61),
	.CK(clk__L2_N4), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[7]  (
	.RN(n54),
	.QN(n78),
	.Q(dataOut[7]),
	.D(n62),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[6]  (
	.RN(n54),
	.QN(n79),
	.Q(dataOut[6]),
	.D(n63),
	.CK(clk__L2_N4), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[5]  (
	.RN(n54),
	.QN(n80),
	.Q(dataOut[5]),
	.D(n64),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[4]  (
	.RN(n54),
	.QN(n81),
	.Q(dataOut[4]),
	.D(n65),
	.CK(clk__L2_N13), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[3]  (
	.RN(n54),
	.QN(n82),
	.Q(dataOut[3]),
	.D(n66),
	.CK(clk__L2_N13), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[2]  (
	.RN(n54),
	.QN(n83),
	.Q(dataOut[2]),
	.D(n67),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[1]  (
	.RN(n54),
	.QN(n84),
	.Q(dataOut[1]),
	.D(n68),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[0]  (
	.RN(n54),
	.QN(n85),
	.Q(dataOut[0]),
	.D(n69),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U2 (
	.ZN(n69),
	.B2(n85),
	.B1(write),
	.A(n101), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U3 (
	.ZN(n101),
	.A2(data[0]),
	.A1(write), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U4 (
	.ZN(n68),
	.B2(n84),
	.B1(write),
	.A(n100), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U5 (
	.ZN(n100),
	.A2(write),
	.A1(data[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U6 (
	.ZN(n67),
	.B2(n83),
	.B1(write),
	.A(n99), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U7 (
	.ZN(n99),
	.A2(write),
	.A1(data[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U8 (
	.ZN(n66),
	.B2(n82),
	.B1(write),
	.A(n98), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U9 (
	.ZN(n98),
	.A2(write),
	.A1(data[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U10 (
	.ZN(n65),
	.B2(n81),
	.B1(write),
	.A(n97), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U11 (
	.ZN(n97),
	.A2(write),
	.A1(data[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U12 (
	.ZN(n64),
	.B2(n80),
	.B1(FE_OFN39_write),
	.A(n96), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U13 (
	.ZN(n96),
	.A2(FE_OFN39_write),
	.A1(data[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U14 (
	.ZN(n63),
	.B2(n79),
	.B1(FE_OFN37_write),
	.A(n95), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U15 (
	.ZN(n95),
	.A2(FE_OFN37_write),
	.A1(data[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U16 (
	.ZN(n62),
	.B2(n78),
	.B1(write),
	.A(n94), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U17 (
	.ZN(n94),
	.A2(write),
	.A1(data[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U18 (
	.ZN(n61),
	.B2(n77),
	.B1(FE_OFN37_write),
	.A(n93), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U19 (
	.ZN(n93),
	.A2(FE_OFN8_write),
	.A1(data[8]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U20 (
	.ZN(n60),
	.B2(n76),
	.B1(write),
	.A(n92), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U21 (
	.ZN(n92),
	.A2(write),
	.A1(data[9]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U22 (
	.ZN(n59),
	.B2(n75),
	.B1(FE_OFN8_write),
	.A(n91), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U23 (
	.ZN(n91),
	.A2(FE_OFN8_write),
	.A1(data[10]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U24 (
	.ZN(n58),
	.B2(n74),
	.B1(FE_OFN37_write),
	.A(n90), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U25 (
	.ZN(n90),
	.A2(FE_OFN37_write),
	.A1(data[11]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U26 (
	.ZN(n57),
	.B2(n73),
	.B1(FE_OFN8_write),
	.A(n89), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U27 (
	.ZN(n89),
	.A2(FE_OFN35_write),
	.A1(data[12]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U28 (
	.ZN(n56),
	.B2(n72),
	.B1(FE_OFN8_write),
	.A(n88), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U29 (
	.ZN(n88),
	.A2(FE_OFN8_write),
	.A1(data[13]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U30 (
	.ZN(n55),
	.B2(n71),
	.B1(FE_OFN35_write),
	.A(n87), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U31 (
	.ZN(n87),
	.A2(FE_OFN35_write),
	.A1(data[14]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U32 (
	.ZN(n54),
	.A(reset), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U33 (
	.ZN(n53),
	.B2(n70),
	.B1(FE_OFN8_write),
	.A(n86), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U34 (
	.ZN(n86),
	.A2(FE_OFN35_write),
	.A1(data[15]), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module SingleReg_3 (
	data, 
	clk, 
	reset, 
	write, 
	dataOut, 
	FE_OFN14_write, 
	FE_OFN9_write, 
	clk__L2_N6, 
	clk__L2_N9, 
	VDD, 
	VSS);
   input [15:0] data;
   input clk;
   input reset;
   input write;
   output [15:0] dataOut;
   input FE_OFN14_write;
   input FE_OFN9_write;
   input clk__L2_N6;
   input clk__L2_N9;
   inout VDD;
   inout VSS;

   // Internal wires
   wire n53;
   wire n54;
   wire n55;
   wire n56;
   wire n57;
   wire n58;
   wire n59;
   wire n60;
   wire n61;
   wire n62;
   wire n63;
   wire n64;
   wire n65;
   wire n66;
   wire n67;
   wire n68;
   wire n69;
   wire n70;
   wire n71;
   wire n72;
   wire n73;
   wire n74;
   wire n75;
   wire n76;
   wire n77;
   wire n78;
   wire n79;
   wire n80;
   wire n81;
   wire n82;
   wire n83;
   wire n84;
   wire n85;
   wire n86;
   wire n87;
   wire n88;
   wire n89;
   wire n90;
   wire n91;
   wire n92;
   wire n93;
   wire n94;
   wire n95;
   wire n96;
   wire n97;
   wire n98;
   wire n99;
   wire n100;
   wire n101;

   // Module instantiations
   DFFR_X1 \Reg_reg[15]  (
	.RN(n54),
	.QN(n70),
	.Q(dataOut[15]),
	.D(n53),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[14]  (
	.RN(n54),
	.QN(n71),
	.Q(dataOut[14]),
	.D(n55),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[13]  (
	.RN(n54),
	.QN(n72),
	.Q(dataOut[13]),
	.D(n56),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[12]  (
	.RN(n54),
	.QN(n73),
	.Q(dataOut[12]),
	.D(n57),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[11]  (
	.RN(n54),
	.QN(n74),
	.Q(dataOut[11]),
	.D(n58),
	.CK(clk__L2_N6), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[10]  (
	.RN(n54),
	.QN(n75),
	.Q(dataOut[10]),
	.D(n59),
	.CK(clk__L2_N6), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[9]  (
	.RN(n54),
	.QN(n76),
	.Q(dataOut[9]),
	.D(n60),
	.CK(clk__L2_N9), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[8]  (
	.RN(n54),
	.QN(n77),
	.Q(dataOut[8]),
	.D(n61),
	.CK(clk__L2_N6), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[7]  (
	.RN(n54),
	.QN(n78),
	.Q(dataOut[7]),
	.D(n62),
	.CK(clk__L2_N9), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[6]  (
	.RN(n54),
	.QN(n79),
	.Q(dataOut[6]),
	.D(n63),
	.CK(clk__L2_N9), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[5]  (
	.RN(n54),
	.QN(n80),
	.Q(dataOut[5]),
	.D(n64),
	.CK(clk__L2_N6), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[4]  (
	.RN(n54),
	.QN(n81),
	.Q(dataOut[4]),
	.D(n65),
	.CK(clk__L2_N9), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[3]  (
	.RN(n54),
	.QN(n82),
	.Q(dataOut[3]),
	.D(n66),
	.CK(clk__L2_N9), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[2]  (
	.RN(n54),
	.QN(n83),
	.Q(dataOut[2]),
	.D(n67),
	.CK(clk__L2_N9), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[1]  (
	.RN(n54),
	.QN(n84),
	.Q(dataOut[1]),
	.D(n68),
	.CK(clk__L2_N9), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[0]  (
	.RN(n54),
	.QN(n85),
	.Q(dataOut[0]),
	.D(n69),
	.CK(clk__L2_N9), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U2 (
	.ZN(n69),
	.B2(n85),
	.B1(FE_OFN14_write),
	.A(n101), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U3 (
	.ZN(n101),
	.A2(data[0]),
	.A1(FE_OFN14_write), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U4 (
	.ZN(n68),
	.B2(n84),
	.B1(FE_OFN14_write),
	.A(n100), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U5 (
	.ZN(n100),
	.A2(FE_OFN14_write),
	.A1(data[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U6 (
	.ZN(n67),
	.B2(n83),
	.B1(FE_OFN14_write),
	.A(n99), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U7 (
	.ZN(n99),
	.A2(FE_OFN14_write),
	.A1(data[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U8 (
	.ZN(n66),
	.B2(n82),
	.B1(FE_OFN14_write),
	.A(n98), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U9 (
	.ZN(n98),
	.A2(FE_OFN14_write),
	.A1(data[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U10 (
	.ZN(n65),
	.B2(n81),
	.B1(FE_OFN14_write),
	.A(n97), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U11 (
	.ZN(n97),
	.A2(FE_OFN14_write),
	.A1(data[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U12 (
	.ZN(n64),
	.B2(n80),
	.B1(FE_OFN14_write),
	.A(n96), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U13 (
	.ZN(n96),
	.A2(FE_OFN14_write),
	.A1(data[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U14 (
	.ZN(n63),
	.B2(n79),
	.B1(FE_OFN14_write),
	.A(n95), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U15 (
	.ZN(n95),
	.A2(FE_OFN14_write),
	.A1(data[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U16 (
	.ZN(n62),
	.B2(n78),
	.B1(FE_OFN14_write),
	.A(n94), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U17 (
	.ZN(n94),
	.A2(FE_OFN14_write),
	.A1(data[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U18 (
	.ZN(n61),
	.B2(n77),
	.B1(FE_OFN14_write),
	.A(n93), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U19 (
	.ZN(n93),
	.A2(FE_OFN14_write),
	.A1(data[8]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U20 (
	.ZN(n60),
	.B2(n76),
	.B1(FE_OFN14_write),
	.A(n92), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U21 (
	.ZN(n92),
	.A2(FE_OFN14_write),
	.A1(data[9]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U22 (
	.ZN(n59),
	.B2(n75),
	.B1(write),
	.A(n91), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U23 (
	.ZN(n91),
	.A2(write),
	.A1(data[10]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U24 (
	.ZN(n58),
	.B2(n74),
	.B1(FE_OFN14_write),
	.A(n90), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U25 (
	.ZN(n90),
	.A2(FE_OFN14_write),
	.A1(data[11]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U26 (
	.ZN(n57),
	.B2(n73),
	.B1(write),
	.A(n89), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U27 (
	.ZN(n89),
	.A2(write),
	.A1(data[12]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U28 (
	.ZN(n56),
	.B2(n72),
	.B1(FE_OFN9_write),
	.A(n88), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U29 (
	.ZN(n88),
	.A2(FE_OFN9_write),
	.A1(data[13]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U30 (
	.ZN(n55),
	.B2(n71),
	.B1(write),
	.A(n87), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U31 (
	.ZN(n87),
	.A2(write),
	.A1(data[14]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U32 (
	.ZN(n54),
	.A(reset), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U33 (
	.ZN(n53),
	.B2(n70),
	.B1(write),
	.A(n86), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U34 (
	.ZN(n86),
	.A2(write),
	.A1(data[15]), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module SingleReg_2 (
	data, 
	clk, 
	reset, 
	write, 
	dataOut, 
	FE_OFN14_write, 
	clk__L2_N6, 
	clk__L2_N9, 
	VDD, 
	VSS);
   input [15:0] data;
   input clk;
   input reset;
   input write;
   output [15:0] dataOut;
   input FE_OFN14_write;
   input clk__L2_N6;
   input clk__L2_N9;
   inout VDD;
   inout VSS;

   // Internal wires
   wire n53;
   wire n54;
   wire n55;
   wire n56;
   wire n57;
   wire n58;
   wire n59;
   wire n60;
   wire n61;
   wire n62;
   wire n63;
   wire n64;
   wire n65;
   wire n66;
   wire n67;
   wire n68;
   wire n69;
   wire n70;
   wire n71;
   wire n72;
   wire n73;
   wire n74;
   wire n75;
   wire n76;
   wire n77;
   wire n78;
   wire n79;
   wire n80;
   wire n81;
   wire n82;
   wire n83;
   wire n84;
   wire n85;
   wire n86;
   wire n87;
   wire n88;
   wire n89;
   wire n90;
   wire n91;
   wire n92;
   wire n93;
   wire n94;
   wire n95;
   wire n96;
   wire n97;
   wire n98;
   wire n99;
   wire n100;
   wire n101;

   // Module instantiations
   DFFR_X1 \Reg_reg[15]  (
	.RN(n54),
	.QN(n70),
	.Q(dataOut[15]),
	.D(n53),
	.CK(clk__L2_N6), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[14]  (
	.RN(n54),
	.QN(n71),
	.Q(dataOut[14]),
	.D(n55),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[13]  (
	.RN(n54),
	.QN(n72),
	.Q(dataOut[13]),
	.D(n56),
	.CK(clk__L2_N6), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[12]  (
	.RN(n54),
	.QN(n73),
	.Q(dataOut[12]),
	.D(n57),
	.CK(clk__L2_N6), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[11]  (
	.RN(n54),
	.QN(n74),
	.Q(dataOut[11]),
	.D(n58),
	.CK(clk__L2_N6), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[10]  (
	.RN(n54),
	.QN(n75),
	.Q(dataOut[10]),
	.D(n59),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[9]  (
	.RN(n54),
	.QN(n76),
	.Q(dataOut[9]),
	.D(n60),
	.CK(clk__L2_N9), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[8]  (
	.RN(n54),
	.QN(n77),
	.Q(dataOut[8]),
	.D(n61),
	.CK(clk__L2_N6), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[7]  (
	.RN(n54),
	.QN(n78),
	.Q(dataOut[7]),
	.D(n62),
	.CK(clk__L2_N9), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[6]  (
	.RN(n54),
	.QN(n79),
	.Q(dataOut[6]),
	.D(n63),
	.CK(clk__L2_N9), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[5]  (
	.RN(n54),
	.QN(n80),
	.Q(dataOut[5]),
	.D(n64),
	.CK(clk__L2_N6), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[4]  (
	.RN(n54),
	.QN(n81),
	.Q(dataOut[4]),
	.D(n65),
	.CK(clk__L2_N9), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[3]  (
	.RN(n54),
	.QN(n82),
	.Q(dataOut[3]),
	.D(n66),
	.CK(clk__L2_N9), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[2]  (
	.RN(n54),
	.QN(n83),
	.Q(dataOut[2]),
	.D(n67),
	.CK(clk__L2_N9), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[1]  (
	.RN(n54),
	.QN(n84),
	.Q(dataOut[1]),
	.D(n68),
	.CK(clk__L2_N9), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[0]  (
	.RN(n54),
	.QN(n85),
	.Q(dataOut[0]),
	.D(n69),
	.CK(clk__L2_N9), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U2 (
	.ZN(n69),
	.B2(n85),
	.B1(FE_OFN14_write),
	.A(n101), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U3 (
	.ZN(n101),
	.A2(data[0]),
	.A1(FE_OFN14_write), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U4 (
	.ZN(n68),
	.B2(n84),
	.B1(FE_OFN14_write),
	.A(n100), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U5 (
	.ZN(n100),
	.A2(FE_OFN14_write),
	.A1(data[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U6 (
	.ZN(n67),
	.B2(n83),
	.B1(FE_OFN14_write),
	.A(n99), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U7 (
	.ZN(n99),
	.A2(FE_OFN14_write),
	.A1(data[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U8 (
	.ZN(n66),
	.B2(n82),
	.B1(FE_OFN14_write),
	.A(n98), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U9 (
	.ZN(n98),
	.A2(FE_OFN14_write),
	.A1(data[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U10 (
	.ZN(n65),
	.B2(n81),
	.B1(FE_OFN14_write),
	.A(n97), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U11 (
	.ZN(n97),
	.A2(FE_OFN14_write),
	.A1(data[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U12 (
	.ZN(n64),
	.B2(n80),
	.B1(FE_OFN14_write),
	.A(n96), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U13 (
	.ZN(n96),
	.A2(FE_OFN14_write),
	.A1(data[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U14 (
	.ZN(n63),
	.B2(n79),
	.B1(FE_OFN14_write),
	.A(n95), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U15 (
	.ZN(n95),
	.A2(FE_OFN14_write),
	.A1(data[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U16 (
	.ZN(n62),
	.B2(n78),
	.B1(FE_OFN14_write),
	.A(n94), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U17 (
	.ZN(n94),
	.A2(FE_OFN14_write),
	.A1(data[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U18 (
	.ZN(n61),
	.B2(n77),
	.B1(FE_OFN14_write),
	.A(n93), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U19 (
	.ZN(n93),
	.A2(FE_OFN14_write),
	.A1(data[8]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U20 (
	.ZN(n60),
	.B2(n76),
	.B1(FE_OFN14_write),
	.A(n92), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U21 (
	.ZN(n92),
	.A2(FE_OFN14_write),
	.A1(data[9]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U22 (
	.ZN(n59),
	.B2(n75),
	.B1(write),
	.A(n91), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U23 (
	.ZN(n91),
	.A2(write),
	.A1(data[10]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U24 (
	.ZN(n58),
	.B2(n74),
	.B1(FE_OFN14_write),
	.A(n90), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U25 (
	.ZN(n90),
	.A2(FE_OFN14_write),
	.A1(data[11]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U26 (
	.ZN(n57),
	.B2(n73),
	.B1(write),
	.A(n89), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U27 (
	.ZN(n89),
	.A2(write),
	.A1(data[12]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U28 (
	.ZN(n56),
	.B2(n72),
	.B1(write),
	.A(n88), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U29 (
	.ZN(n88),
	.A2(write),
	.A1(data[13]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U30 (
	.ZN(n55),
	.B2(n71),
	.B1(write),
	.A(n87), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U31 (
	.ZN(n87),
	.A2(write),
	.A1(data[14]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U32 (
	.ZN(n54),
	.A(reset), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U33 (
	.ZN(n53),
	.B2(n70),
	.B1(write),
	.A(n86), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U34 (
	.ZN(n86),
	.A2(write),
	.A1(data[15]), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module SingleReg_1 (
	data, 
	clk, 
	reset, 
	write, 
	dataOut, 
	FE_OFN13_write, 
	FE_OFN14_write, 
	FE_OFN57_write, 
	FE_OFN58_write, 
	FE_OFN59_write, 
	clk__L2_N9, 
	VDD, 
	VSS);
   input [15:0] data;
   input clk;
   input reset;
   input write;
   output [15:0] dataOut;
   input FE_OFN13_write;
   input FE_OFN14_write;
   input FE_OFN57_write;
   input FE_OFN58_write;
   input FE_OFN59_write;
   input clk__L2_N9;
   inout VDD;
   inout VSS;

   // Internal wires
   wire n53;
   wire n54;
   wire n55;
   wire n56;
   wire n57;
   wire n58;
   wire n59;
   wire n60;
   wire n61;
   wire n62;
   wire n63;
   wire n64;
   wire n65;
   wire n66;
   wire n67;
   wire n68;
   wire n69;
   wire n70;
   wire n71;
   wire n72;
   wire n73;
   wire n74;
   wire n75;
   wire n76;
   wire n77;
   wire n78;
   wire n79;
   wire n80;
   wire n81;
   wire n82;
   wire n83;
   wire n84;
   wire n85;
   wire n86;
   wire n87;
   wire n88;
   wire n89;
   wire n90;
   wire n91;
   wire n92;
   wire n93;
   wire n94;
   wire n95;
   wire n96;
   wire n97;
   wire n98;
   wire n99;
   wire n100;
   wire n101;

   // Module instantiations
   DFFR_X1 \Reg_reg[15]  (
	.RN(n54),
	.QN(n70),
	.Q(dataOut[15]),
	.D(n53),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[14]  (
	.RN(n54),
	.QN(n71),
	.Q(dataOut[14]),
	.D(n55),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[13]  (
	.RN(n54),
	.QN(n72),
	.Q(dataOut[13]),
	.D(n56),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[12]  (
	.RN(n54),
	.QN(n73),
	.Q(dataOut[12]),
	.D(n57),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[11]  (
	.RN(n54),
	.QN(n74),
	.Q(dataOut[11]),
	.D(n58),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[10]  (
	.RN(n54),
	.QN(n75),
	.Q(dataOut[10]),
	.D(n59),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[9]  (
	.RN(n54),
	.QN(n76),
	.Q(dataOut[9]),
	.D(n60),
	.CK(clk__L2_N9), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[8]  (
	.RN(n54),
	.QN(n77),
	.Q(dataOut[8]),
	.D(n61),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[7]  (
	.RN(n54),
	.QN(n78),
	.Q(dataOut[7]),
	.D(n62),
	.CK(clk__L2_N9), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[6]  (
	.RN(n54),
	.QN(n79),
	.Q(dataOut[6]),
	.D(n63),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[5]  (
	.RN(n54),
	.QN(n80),
	.Q(dataOut[5]),
	.D(n64),
	.CK(clk__L2_N9), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[4]  (
	.RN(n54),
	.QN(n81),
	.Q(dataOut[4]),
	.D(n65),
	.CK(clk__L2_N9), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[3]  (
	.RN(n54),
	.QN(n82),
	.Q(dataOut[3]),
	.D(n66),
	.CK(clk__L2_N9), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[2]  (
	.RN(n54),
	.QN(n83),
	.Q(dataOut[2]),
	.D(n67),
	.CK(clk__L2_N9), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[1]  (
	.RN(n54),
	.QN(n84),
	.Q(dataOut[1]),
	.D(n68),
	.CK(clk__L2_N9), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[0]  (
	.RN(n54),
	.QN(n85),
	.Q(dataOut[0]),
	.D(n69),
	.CK(clk__L2_N9), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U2 (
	.ZN(n69),
	.B2(n85),
	.B1(write),
	.A(n101), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U3 (
	.ZN(n101),
	.A2(data[0]),
	.A1(write), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U4 (
	.ZN(n68),
	.B2(n84),
	.B1(write),
	.A(n100), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U5 (
	.ZN(n100),
	.A2(write),
	.A1(data[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U6 (
	.ZN(n67),
	.B2(n83),
	.B1(FE_OFN14_write),
	.A(n99), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U7 (
	.ZN(n99),
	.A2(FE_OFN14_write),
	.A1(data[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U8 (
	.ZN(n66),
	.B2(n82),
	.B1(FE_OFN14_write),
	.A(n98), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U9 (
	.ZN(n98),
	.A2(write),
	.A1(data[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U10 (
	.ZN(n65),
	.B2(n81),
	.B1(FE_OFN58_write),
	.A(n97), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U11 (
	.ZN(n97),
	.A2(FE_OFN58_write),
	.A1(data[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U12 (
	.ZN(n64),
	.B2(n80),
	.B1(FE_OFN13_write),
	.A(n96), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U13 (
	.ZN(n96),
	.A2(FE_OFN14_write),
	.A1(data[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U14 (
	.ZN(n63),
	.B2(n79),
	.B1(FE_OFN59_write),
	.A(n95), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U15 (
	.ZN(n95),
	.A2(FE_OFN57_write),
	.A1(data[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U16 (
	.ZN(n62),
	.B2(n78),
	.B1(write),
	.A(n94), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U17 (
	.ZN(n94),
	.A2(write),
	.A1(data[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U18 (
	.ZN(n61),
	.B2(n77),
	.B1(FE_OFN59_write),
	.A(n93), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U19 (
	.ZN(n93),
	.A2(FE_OFN59_write),
	.A1(data[8]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U20 (
	.ZN(n60),
	.B2(n76),
	.B1(FE_OFN58_write),
	.A(n92), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U21 (
	.ZN(n92),
	.A2(FE_OFN58_write),
	.A1(data[9]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U22 (
	.ZN(n59),
	.B2(n75),
	.B1(FE_OFN59_write),
	.A(n91), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U23 (
	.ZN(n91),
	.A2(FE_OFN59_write),
	.A1(data[10]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U24 (
	.ZN(n58),
	.B2(n74),
	.B1(FE_OFN13_write),
	.A(n90), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U25 (
	.ZN(n90),
	.A2(FE_OFN13_write),
	.A1(data[11]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U26 (
	.ZN(n57),
	.B2(n73),
	.B1(FE_OFN57_write),
	.A(n89), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U27 (
	.ZN(n89),
	.A2(FE_OFN57_write),
	.A1(data[12]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U28 (
	.ZN(n56),
	.B2(n72),
	.B1(FE_OFN59_write),
	.A(n88), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U29 (
	.ZN(n88),
	.A2(FE_OFN59_write),
	.A1(data[13]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U30 (
	.ZN(n55),
	.B2(n71),
	.B1(FE_OFN59_write),
	.A(n87), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U31 (
	.ZN(n87),
	.A2(FE_OFN59_write),
	.A1(data[14]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U32 (
	.ZN(n54),
	.A(reset), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U33 (
	.ZN(n53),
	.B2(n70),
	.B1(FE_OFN57_write),
	.A(n86), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U34 (
	.ZN(n86),
	.A2(FE_OFN57_write),
	.A1(data[15]), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module SingleReg_0 (
	data, 
	clk, 
	reset, 
	write, 
	dataOut, 
	FE_OFN13_write, 
	FE_OFN14_write, 
	FE_OFN9_write, 
	FE_OFN57_write, 
	FE_OFN58_write, 
	FE_OFN59_write, 
	clk__L2_N6, 
	clk__L2_N9, 
	VDD, 
	VSS);
   input [15:0] data;
   input clk;
   input reset;
   input write;
   output [15:0] dataOut;
   input FE_OFN13_write;
   input FE_OFN14_write;
   input FE_OFN9_write;
   input FE_OFN57_write;
   input FE_OFN58_write;
   input FE_OFN59_write;
   input clk__L2_N6;
   input clk__L2_N9;
   inout VDD;
   inout VSS;

   // Internal wires
   wire n53;
   wire n54;
   wire n55;
   wire n56;
   wire n57;
   wire n58;
   wire n59;
   wire n60;
   wire n61;
   wire n62;
   wire n63;
   wire n64;
   wire n65;
   wire n66;
   wire n67;
   wire n68;
   wire n69;
   wire n70;
   wire n71;
   wire n72;
   wire n73;
   wire n74;
   wire n75;
   wire n76;
   wire n77;
   wire n78;
   wire n79;
   wire n80;
   wire n81;
   wire n82;
   wire n83;
   wire n84;
   wire n85;
   wire n86;
   wire n87;
   wire n88;
   wire n89;
   wire n90;
   wire n91;
   wire n92;
   wire n93;
   wire n94;
   wire n95;
   wire n96;
   wire n97;
   wire n98;
   wire n99;
   wire n100;
   wire n101;

   // Module instantiations
   DFFR_X1 \Reg_reg[15]  (
	.RN(n54),
	.QN(n70),
	.Q(dataOut[15]),
	.D(n53),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[14]  (
	.RN(n54),
	.QN(n71),
	.Q(dataOut[14]),
	.D(n55),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[13]  (
	.RN(n54),
	.QN(n72),
	.Q(dataOut[13]),
	.D(n56),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[12]  (
	.RN(n54),
	.QN(n73),
	.Q(dataOut[12]),
	.D(n57),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[11]  (
	.RN(n54),
	.QN(n74),
	.Q(dataOut[11]),
	.D(n58),
	.CK(clk__L2_N6), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[10]  (
	.RN(n54),
	.QN(n75),
	.Q(dataOut[10]),
	.D(n59),
	.CK(clk__L2_N6), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[9]  (
	.RN(n54),
	.QN(n76),
	.Q(dataOut[9]),
	.D(n60),
	.CK(clk__L2_N9), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[8]  (
	.RN(n54),
	.QN(n77),
	.Q(dataOut[8]),
	.D(n61),
	.CK(clk__L2_N6), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[7]  (
	.RN(n54),
	.QN(n78),
	.Q(dataOut[7]),
	.D(n62),
	.CK(clk__L2_N9), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[6]  (
	.RN(n54),
	.QN(n79),
	.Q(dataOut[6]),
	.D(n63),
	.CK(clk__L2_N6), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[5]  (
	.RN(n54),
	.QN(n80),
	.Q(dataOut[5]),
	.D(n64),
	.CK(clk__L2_N9), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[4]  (
	.RN(n54),
	.QN(n81),
	.Q(dataOut[4]),
	.D(n65),
	.CK(clk__L2_N9), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[3]  (
	.RN(n54),
	.QN(n82),
	.Q(dataOut[3]),
	.D(n66),
	.CK(clk__L2_N9), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[2]  (
	.RN(n54),
	.QN(n83),
	.Q(dataOut[2]),
	.D(n67),
	.CK(clk__L2_N9), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[1]  (
	.RN(n54),
	.QN(n84),
	.Q(dataOut[1]),
	.D(n68),
	.CK(clk__L2_N9), 
	.VDD(VDD), 
	.VSS(VSS));
   DFFR_X1 \Reg_reg[0]  (
	.RN(n54),
	.QN(n85),
	.Q(dataOut[0]),
	.D(n69),
	.CK(clk__L2_N9), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U2 (
	.ZN(n69),
	.B2(n85),
	.B1(write),
	.A(n101), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U3 (
	.ZN(n101),
	.A2(data[0]),
	.A1(write), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U4 (
	.ZN(n68),
	.B2(n84),
	.B1(write),
	.A(n100), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U5 (
	.ZN(n100),
	.A2(write),
	.A1(data[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U6 (
	.ZN(n67),
	.B2(n83),
	.B1(FE_OFN14_write),
	.A(n99), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U7 (
	.ZN(n99),
	.A2(FE_OFN14_write),
	.A1(data[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U8 (
	.ZN(n66),
	.B2(n82),
	.B1(FE_OFN14_write),
	.A(n98), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U9 (
	.ZN(n98),
	.A2(FE_OFN14_write),
	.A1(data[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U10 (
	.ZN(n65),
	.B2(n81),
	.B1(FE_OFN14_write),
	.A(n97), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U11 (
	.ZN(n97),
	.A2(FE_OFN58_write),
	.A1(data[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U12 (
	.ZN(n64),
	.B2(n80),
	.B1(FE_OFN14_write),
	.A(n96), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U13 (
	.ZN(n96),
	.A2(FE_OFN14_write),
	.A1(data[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U14 (
	.ZN(n63),
	.B2(n79),
	.B1(FE_OFN13_write),
	.A(n95), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U15 (
	.ZN(n95),
	.A2(FE_OFN13_write),
	.A1(data[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U16 (
	.ZN(n62),
	.B2(n78),
	.B1(write),
	.A(n94), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U17 (
	.ZN(n94),
	.A2(write),
	.A1(data[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U18 (
	.ZN(n61),
	.B2(n77),
	.B1(FE_OFN57_write),
	.A(n93), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U19 (
	.ZN(n93),
	.A2(FE_OFN57_write),
	.A1(data[8]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U20 (
	.ZN(n60),
	.B2(n76),
	.B1(write),
	.A(n92), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U21 (
	.ZN(n92),
	.A2(write),
	.A1(data[9]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U22 (
	.ZN(n59),
	.B2(n75),
	.B1(FE_OFN59_write),
	.A(n91), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U23 (
	.ZN(n91),
	.A2(FE_OFN59_write),
	.A1(data[10]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U24 (
	.ZN(n58),
	.B2(n74),
	.B1(FE_OFN59_write),
	.A(n90), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U25 (
	.ZN(n90),
	.A2(FE_OFN59_write),
	.A1(data[11]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U26 (
	.ZN(n57),
	.B2(n73),
	.B1(FE_OFN9_write),
	.A(n89), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U27 (
	.ZN(n89),
	.A2(FE_OFN9_write),
	.A1(data[12]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U28 (
	.ZN(n56),
	.B2(n72),
	.B1(FE_OFN59_write),
	.A(n88), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U29 (
	.ZN(n88),
	.A2(FE_OFN59_write),
	.A1(data[13]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U30 (
	.ZN(n55),
	.B2(n71),
	.B1(FE_OFN59_write),
	.A(n87), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U31 (
	.ZN(n87),
	.A2(FE_OFN59_write),
	.A1(data[14]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X2 U32 (
	.ZN(n54),
	.A(reset), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21_X1 U33 (
	.ZN(n53),
	.B2(n70),
	.B1(FE_OFN59_write),
	.A(n86), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U34 (
	.ZN(n86),
	.A2(FE_OFN59_write),
	.A1(data[15]), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module RegFile (
	addressA, 
	addressB, 
	dataIn, 
	addressIn, 
	clk, 
	reset, 
	write, 
	outA, 
	outB, 
	VDD, 
	VSS);
   input [4:0] addressA;
   input [4:0] addressB;
   input [15:0] dataIn;
   input [4:0] addressIn;
   input clk;
   input reset;
   input write;
   output [15:0] outA;
   output [15:0] outB;
   inout VDD;
   inout VSS;

   // Internal wires
   wire clk__L2_N13;
   wire clk__L2_N12;
   wire clk__L2_N11;
   wire clk__L2_N10;
   wire clk__L2_N9;
   wire clk__L2_N8;
   wire clk__L2_N7;
   wire clk__L2_N6;
   wire clk__L2_N5;
   wire clk__L2_N4;
   wire clk__L2_N3;
   wire clk__L2_N2;
   wire clk__L2_N1;
   wire clk__L2_N0;
   wire clk__L1_N0;
   wire FE_UNCONNECTED_0;
   wire FE_OFN75_n569;
   wire FE_OFN74_n568;
   wire FE_OFN73_n574;
   wire FE_OFN72_n573;
   wire FE_OFN71_n603;
   wire FE_OFN70_n602;
   wire FE_OFN69_n608;
   wire FE_OFN68_n607;
   wire FE_OFN67_n579;
   wire FE_OFN66_n578;
   wire FE_OFN65_n584;
   wire FE_OFN64_n583;
   wire FE_OFN63_n593;
   wire FE_OFN62_n592;
   wire FE_OFN61_n598;
   wire FE_OFN60_n597;
   wire FE_OFN59_write;
   wire FE_OFN58_write;
   wire FE_OFN57_write;
   wire FE_OFN56_write;
   wire FE_OFN55_write;
   wire FE_OFN54_write;
   wire FE_OFN53_write;
   wire FE_OFN51_write;
   wire FE_OFN50_write;
   wire FE_OFN49_write;
   wire FE_OFN48_write;
   wire FE_OFN47_write;
   wire FE_OFN46_write;
   wire FE_OFN45_write;
   wire FE_OFN44_write;
   wire FE_OFN43_write;
   wire FE_OFN42_write;
   wire FE_OFN41_write;
   wire FE_OFN40_write;
   wire FE_OFN39_write;
   wire FE_OFN38_write;
   wire FE_OFN35_write;
   wire FE_OFN34_write;
   wire FE_OFN32_write;
   wire FE_OFN31_write;
   wire FE_OFN30_write;
   wire FE_OFN29_write;
   wire FE_OFN28_write;
   wire FE_OFN26_write;
   wire FE_OFN25_write;
   wire FE_OFN24_write;
   wire FE_OFN23_write;
   wire FE_OFN22_write;
   wire FE_OFN21_write;
   wire FE_OFN20_write;
   wire FE_OFN18_write;
   wire FE_OFN17_write;
   wire FE_OFN16_write;
   wire FE_OFN15_write;
   wire \regOut[0][15] ;
   wire \regOut[0][14] ;
   wire \regOut[0][13] ;
   wire \regOut[0][12] ;
   wire \regOut[0][11] ;
   wire \regOut[0][10] ;
   wire \regOut[0][9] ;
   wire \regOut[0][8] ;
   wire \regOut[0][7] ;
   wire \regOut[0][6] ;
   wire \regOut[0][5] ;
   wire \regOut[0][4] ;
   wire \regOut[0][3] ;
   wire \regOut[0][2] ;
   wire \regOut[0][1] ;
   wire \regOut[0][0] ;
   wire \regOut[1][15] ;
   wire \regOut[1][14] ;
   wire \regOut[1][13] ;
   wire \regOut[1][12] ;
   wire \regOut[1][11] ;
   wire \regOut[1][10] ;
   wire \regOut[1][9] ;
   wire \regOut[1][8] ;
   wire \regOut[1][7] ;
   wire \regOut[1][6] ;
   wire \regOut[1][5] ;
   wire \regOut[1][4] ;
   wire \regOut[1][3] ;
   wire \regOut[1][2] ;
   wire \regOut[1][1] ;
   wire \regOut[1][0] ;
   wire \regOut[2][15] ;
   wire \regOut[2][14] ;
   wire \regOut[2][13] ;
   wire \regOut[2][12] ;
   wire \regOut[2][11] ;
   wire \regOut[2][10] ;
   wire \regOut[2][9] ;
   wire \regOut[2][8] ;
   wire \regOut[2][7] ;
   wire \regOut[2][6] ;
   wire \regOut[2][5] ;
   wire \regOut[2][4] ;
   wire \regOut[2][3] ;
   wire \regOut[2][2] ;
   wire \regOut[2][1] ;
   wire \regOut[2][0] ;
   wire \regOut[3][15] ;
   wire \regOut[3][14] ;
   wire \regOut[3][13] ;
   wire \regOut[3][12] ;
   wire \regOut[3][11] ;
   wire \regOut[3][10] ;
   wire \regOut[3][9] ;
   wire \regOut[3][8] ;
   wire \regOut[3][7] ;
   wire \regOut[3][6] ;
   wire \regOut[3][5] ;
   wire \regOut[3][4] ;
   wire \regOut[3][3] ;
   wire \regOut[3][2] ;
   wire \regOut[3][1] ;
   wire \regOut[3][0] ;
   wire \regOut[4][15] ;
   wire \regOut[4][14] ;
   wire \regOut[4][13] ;
   wire \regOut[4][12] ;
   wire \regOut[4][11] ;
   wire \regOut[4][10] ;
   wire \regOut[4][9] ;
   wire \regOut[4][8] ;
   wire \regOut[4][7] ;
   wire \regOut[4][6] ;
   wire \regOut[4][5] ;
   wire \regOut[4][4] ;
   wire \regOut[4][3] ;
   wire \regOut[4][2] ;
   wire \regOut[4][1] ;
   wire \regOut[4][0] ;
   wire \regOut[5][15] ;
   wire \regOut[5][14] ;
   wire \regOut[5][13] ;
   wire \regOut[5][12] ;
   wire \regOut[5][11] ;
   wire \regOut[5][10] ;
   wire \regOut[5][9] ;
   wire \regOut[5][8] ;
   wire \regOut[5][7] ;
   wire \regOut[5][6] ;
   wire \regOut[5][5] ;
   wire \regOut[5][4] ;
   wire \regOut[5][3] ;
   wire \regOut[5][2] ;
   wire \regOut[5][1] ;
   wire \regOut[5][0] ;
   wire \regOut[6][15] ;
   wire \regOut[6][14] ;
   wire \regOut[6][13] ;
   wire \regOut[6][12] ;
   wire \regOut[6][11] ;
   wire \regOut[6][10] ;
   wire \regOut[6][9] ;
   wire \regOut[6][8] ;
   wire \regOut[6][7] ;
   wire \regOut[6][6] ;
   wire \regOut[6][5] ;
   wire \regOut[6][4] ;
   wire \regOut[6][3] ;
   wire \regOut[6][2] ;
   wire \regOut[6][1] ;
   wire \regOut[6][0] ;
   wire \regOut[7][15] ;
   wire \regOut[7][14] ;
   wire \regOut[7][13] ;
   wire \regOut[7][12] ;
   wire \regOut[7][11] ;
   wire \regOut[7][10] ;
   wire \regOut[7][9] ;
   wire \regOut[7][8] ;
   wire \regOut[7][7] ;
   wire \regOut[7][6] ;
   wire \regOut[7][5] ;
   wire \regOut[7][4] ;
   wire \regOut[7][3] ;
   wire \regOut[7][2] ;
   wire \regOut[7][1] ;
   wire \regOut[7][0] ;
   wire \regOut[8][15] ;
   wire \regOut[8][14] ;
   wire \regOut[8][13] ;
   wire \regOut[8][12] ;
   wire \regOut[8][11] ;
   wire \regOut[8][10] ;
   wire \regOut[8][9] ;
   wire \regOut[8][8] ;
   wire \regOut[8][7] ;
   wire \regOut[8][6] ;
   wire \regOut[8][5] ;
   wire \regOut[8][4] ;
   wire \regOut[8][3] ;
   wire \regOut[8][2] ;
   wire \regOut[8][1] ;
   wire \regOut[8][0] ;
   wire \regOut[9][15] ;
   wire \regOut[9][14] ;
   wire \regOut[9][13] ;
   wire \regOut[9][12] ;
   wire \regOut[9][11] ;
   wire \regOut[9][10] ;
   wire \regOut[9][9] ;
   wire \regOut[9][8] ;
   wire \regOut[9][7] ;
   wire \regOut[9][6] ;
   wire \regOut[9][5] ;
   wire \regOut[9][4] ;
   wire \regOut[9][3] ;
   wire \regOut[9][2] ;
   wire \regOut[9][1] ;
   wire \regOut[9][0] ;
   wire \regOut[10][15] ;
   wire \regOut[10][14] ;
   wire \regOut[10][13] ;
   wire \regOut[10][12] ;
   wire \regOut[10][11] ;
   wire \regOut[10][10] ;
   wire \regOut[10][9] ;
   wire \regOut[10][8] ;
   wire \regOut[10][7] ;
   wire \regOut[10][6] ;
   wire \regOut[10][5] ;
   wire \regOut[10][4] ;
   wire \regOut[10][3] ;
   wire \regOut[10][2] ;
   wire \regOut[10][1] ;
   wire \regOut[10][0] ;
   wire \regOut[11][15] ;
   wire \regOut[11][14] ;
   wire \regOut[11][13] ;
   wire \regOut[11][12] ;
   wire \regOut[11][11] ;
   wire \regOut[11][10] ;
   wire \regOut[11][9] ;
   wire \regOut[11][8] ;
   wire \regOut[11][7] ;
   wire \regOut[11][6] ;
   wire \regOut[11][5] ;
   wire \regOut[11][4] ;
   wire \regOut[11][3] ;
   wire \regOut[11][2] ;
   wire \regOut[11][1] ;
   wire \regOut[11][0] ;
   wire \regOut[12][15] ;
   wire \regOut[12][14] ;
   wire \regOut[12][13] ;
   wire \regOut[12][12] ;
   wire \regOut[12][11] ;
   wire \regOut[12][10] ;
   wire \regOut[12][9] ;
   wire \regOut[12][8] ;
   wire \regOut[12][7] ;
   wire \regOut[12][6] ;
   wire \regOut[12][5] ;
   wire \regOut[12][4] ;
   wire \regOut[12][3] ;
   wire \regOut[12][2] ;
   wire \regOut[12][1] ;
   wire \regOut[12][0] ;
   wire \regOut[13][15] ;
   wire \regOut[13][14] ;
   wire \regOut[13][13] ;
   wire \regOut[13][12] ;
   wire \regOut[13][11] ;
   wire \regOut[13][10] ;
   wire \regOut[13][9] ;
   wire \regOut[13][8] ;
   wire \regOut[13][7] ;
   wire \regOut[13][6] ;
   wire \regOut[13][5] ;
   wire \regOut[13][4] ;
   wire \regOut[13][3] ;
   wire \regOut[13][2] ;
   wire \regOut[13][1] ;
   wire \regOut[13][0] ;
   wire \regOut[14][15] ;
   wire \regOut[14][14] ;
   wire \regOut[14][13] ;
   wire \regOut[14][12] ;
   wire \regOut[14][11] ;
   wire \regOut[14][10] ;
   wire \regOut[14][9] ;
   wire \regOut[14][8] ;
   wire \regOut[14][7] ;
   wire \regOut[14][6] ;
   wire \regOut[14][5] ;
   wire \regOut[14][4] ;
   wire \regOut[14][3] ;
   wire \regOut[14][2] ;
   wire \regOut[14][1] ;
   wire \regOut[14][0] ;
   wire \regOut[15][15] ;
   wire \regOut[15][14] ;
   wire \regOut[15][13] ;
   wire \regOut[15][12] ;
   wire \regOut[15][11] ;
   wire \regOut[15][10] ;
   wire \regOut[15][9] ;
   wire \regOut[15][8] ;
   wire \regOut[15][7] ;
   wire \regOut[15][6] ;
   wire \regOut[15][5] ;
   wire \regOut[15][4] ;
   wire \regOut[15][3] ;
   wire \regOut[15][2] ;
   wire \regOut[15][1] ;
   wire \regOut[15][0] ;
   wire \regOut[16][15] ;
   wire \regOut[16][14] ;
   wire \regOut[16][13] ;
   wire \regOut[16][12] ;
   wire \regOut[16][11] ;
   wire \regOut[16][10] ;
   wire \regOut[16][9] ;
   wire \regOut[16][8] ;
   wire \regOut[16][7] ;
   wire \regOut[16][6] ;
   wire \regOut[16][5] ;
   wire \regOut[16][4] ;
   wire \regOut[16][3] ;
   wire \regOut[16][2] ;
   wire \regOut[16][1] ;
   wire \regOut[16][0] ;
   wire \regOut[17][15] ;
   wire \regOut[17][14] ;
   wire \regOut[17][13] ;
   wire \regOut[17][12] ;
   wire \regOut[17][11] ;
   wire \regOut[17][10] ;
   wire \regOut[17][9] ;
   wire \regOut[17][8] ;
   wire \regOut[17][7] ;
   wire \regOut[17][6] ;
   wire \regOut[17][5] ;
   wire \regOut[17][4] ;
   wire \regOut[17][3] ;
   wire \regOut[17][2] ;
   wire \regOut[17][1] ;
   wire \regOut[17][0] ;
   wire \regOut[18][15] ;
   wire \regOut[18][14] ;
   wire \regOut[18][13] ;
   wire \regOut[18][12] ;
   wire \regOut[18][11] ;
   wire \regOut[18][10] ;
   wire \regOut[18][9] ;
   wire \regOut[18][8] ;
   wire \regOut[18][7] ;
   wire \regOut[18][6] ;
   wire \regOut[18][5] ;
   wire \regOut[18][4] ;
   wire \regOut[18][3] ;
   wire \regOut[18][2] ;
   wire \regOut[18][1] ;
   wire \regOut[18][0] ;
   wire \regOut[19][15] ;
   wire \regOut[19][14] ;
   wire \regOut[19][13] ;
   wire \regOut[19][12] ;
   wire \regOut[19][11] ;
   wire \regOut[19][10] ;
   wire \regOut[19][9] ;
   wire \regOut[19][8] ;
   wire \regOut[19][7] ;
   wire \regOut[19][6] ;
   wire \regOut[19][5] ;
   wire \regOut[19][4] ;
   wire \regOut[19][3] ;
   wire \regOut[19][2] ;
   wire \regOut[19][1] ;
   wire \regOut[19][0] ;
   wire \regOut[20][15] ;
   wire \regOut[20][14] ;
   wire \regOut[20][13] ;
   wire \regOut[20][12] ;
   wire \regOut[20][11] ;
   wire \regOut[20][10] ;
   wire \regOut[20][9] ;
   wire \regOut[20][8] ;
   wire \regOut[20][7] ;
   wire \regOut[20][6] ;
   wire \regOut[20][5] ;
   wire \regOut[20][4] ;
   wire \regOut[20][3] ;
   wire \regOut[20][2] ;
   wire \regOut[20][1] ;
   wire \regOut[20][0] ;
   wire \regOut[21][15] ;
   wire \regOut[21][14] ;
   wire \regOut[21][13] ;
   wire \regOut[21][12] ;
   wire \regOut[21][11] ;
   wire \regOut[21][10] ;
   wire \regOut[21][9] ;
   wire \regOut[21][8] ;
   wire \regOut[21][7] ;
   wire \regOut[21][6] ;
   wire \regOut[21][5] ;
   wire \regOut[21][4] ;
   wire \regOut[21][3] ;
   wire \regOut[21][2] ;
   wire \regOut[21][1] ;
   wire \regOut[21][0] ;
   wire \regOut[22][15] ;
   wire \regOut[22][14] ;
   wire \regOut[22][13] ;
   wire \regOut[22][12] ;
   wire \regOut[22][11] ;
   wire \regOut[22][10] ;
   wire \regOut[22][9] ;
   wire \regOut[22][8] ;
   wire \regOut[22][7] ;
   wire \regOut[22][6] ;
   wire \regOut[22][5] ;
   wire \regOut[22][4] ;
   wire \regOut[22][3] ;
   wire \regOut[22][2] ;
   wire \regOut[22][1] ;
   wire \regOut[22][0] ;
   wire \regOut[23][15] ;
   wire \regOut[23][14] ;
   wire \regOut[23][13] ;
   wire \regOut[23][12] ;
   wire \regOut[23][11] ;
   wire \regOut[23][10] ;
   wire \regOut[23][9] ;
   wire \regOut[23][8] ;
   wire \regOut[23][7] ;
   wire \regOut[23][6] ;
   wire \regOut[23][5] ;
   wire \regOut[23][4] ;
   wire \regOut[23][3] ;
   wire \regOut[23][2] ;
   wire \regOut[23][1] ;
   wire \regOut[23][0] ;
   wire \regOut[24][15] ;
   wire \regOut[24][14] ;
   wire \regOut[24][13] ;
   wire \regOut[24][12] ;
   wire \regOut[24][11] ;
   wire \regOut[24][10] ;
   wire \regOut[24][9] ;
   wire \regOut[24][8] ;
   wire \regOut[24][7] ;
   wire \regOut[24][6] ;
   wire \regOut[24][5] ;
   wire \regOut[24][4] ;
   wire \regOut[24][3] ;
   wire \regOut[24][2] ;
   wire \regOut[24][1] ;
   wire \regOut[24][0] ;
   wire \regOut[25][15] ;
   wire \regOut[25][14] ;
   wire \regOut[25][13] ;
   wire \regOut[25][12] ;
   wire \regOut[25][11] ;
   wire \regOut[25][10] ;
   wire \regOut[25][9] ;
   wire \regOut[25][8] ;
   wire \regOut[25][7] ;
   wire \regOut[25][6] ;
   wire \regOut[25][5] ;
   wire \regOut[25][4] ;
   wire \regOut[25][3] ;
   wire \regOut[25][2] ;
   wire \regOut[25][1] ;
   wire \regOut[25][0] ;
   wire \regOut[26][15] ;
   wire \regOut[26][14] ;
   wire \regOut[26][13] ;
   wire \regOut[26][12] ;
   wire \regOut[26][11] ;
   wire \regOut[26][10] ;
   wire \regOut[26][9] ;
   wire \regOut[26][8] ;
   wire \regOut[26][7] ;
   wire \regOut[26][6] ;
   wire \regOut[26][5] ;
   wire \regOut[26][4] ;
   wire \regOut[26][3] ;
   wire \regOut[26][2] ;
   wire \regOut[26][1] ;
   wire \regOut[26][0] ;
   wire \regOut[27][15] ;
   wire \regOut[27][14] ;
   wire \regOut[27][13] ;
   wire \regOut[27][12] ;
   wire \regOut[27][11] ;
   wire \regOut[27][10] ;
   wire \regOut[27][9] ;
   wire \regOut[27][8] ;
   wire \regOut[27][7] ;
   wire \regOut[27][6] ;
   wire \regOut[27][5] ;
   wire \regOut[27][4] ;
   wire \regOut[27][3] ;
   wire \regOut[27][2] ;
   wire \regOut[27][1] ;
   wire \regOut[27][0] ;
   wire \regOut[28][15] ;
   wire \regOut[28][14] ;
   wire \regOut[28][13] ;
   wire \regOut[28][12] ;
   wire \regOut[28][11] ;
   wire \regOut[28][10] ;
   wire \regOut[28][9] ;
   wire \regOut[28][8] ;
   wire \regOut[28][7] ;
   wire \regOut[28][6] ;
   wire \regOut[28][5] ;
   wire \regOut[28][4] ;
   wire \regOut[28][3] ;
   wire \regOut[28][2] ;
   wire \regOut[28][1] ;
   wire \regOut[28][0] ;
   wire \regOut[29][15] ;
   wire \regOut[29][14] ;
   wire \regOut[29][13] ;
   wire \regOut[29][12] ;
   wire \regOut[29][11] ;
   wire \regOut[29][10] ;
   wire \regOut[29][9] ;
   wire \regOut[29][8] ;
   wire \regOut[29][7] ;
   wire \regOut[29][6] ;
   wire \regOut[29][5] ;
   wire \regOut[29][4] ;
   wire \regOut[29][3] ;
   wire \regOut[29][2] ;
   wire \regOut[29][1] ;
   wire \regOut[29][0] ;
   wire \regOut[30][15] ;
   wire \regOut[30][14] ;
   wire \regOut[30][13] ;
   wire \regOut[30][12] ;
   wire \regOut[30][11] ;
   wire \regOut[30][10] ;
   wire \regOut[30][9] ;
   wire \regOut[30][8] ;
   wire \regOut[30][7] ;
   wire \regOut[30][6] ;
   wire \regOut[30][5] ;
   wire \regOut[30][4] ;
   wire \regOut[30][3] ;
   wire \regOut[30][2] ;
   wire \regOut[30][1] ;
   wire \regOut[30][0] ;
   wire \regOut[31][15] ;
   wire \regOut[31][14] ;
   wire \regOut[31][13] ;
   wire \regOut[31][12] ;
   wire \regOut[31][11] ;
   wire \regOut[31][10] ;
   wire \regOut[31][9] ;
   wire \regOut[31][8] ;
   wire \regOut[31][7] ;
   wire \regOut[31][6] ;
   wire \regOut[31][5] ;
   wire \regOut[31][4] ;
   wire \regOut[31][3] ;
   wire \regOut[31][2] ;
   wire \regOut[31][1] ;
   wire \regOut[31][0] ;
   wire \regIn[0][15] ;
   wire \regIn[0][14] ;
   wire \regIn[0][13] ;
   wire \regIn[0][12] ;
   wire \regIn[0][11] ;
   wire \regIn[0][10] ;
   wire \regIn[0][9] ;
   wire \regIn[0][8] ;
   wire \regIn[0][7] ;
   wire \regIn[0][6] ;
   wire \regIn[0][5] ;
   wire \regIn[0][4] ;
   wire \regIn[0][3] ;
   wire \regIn[0][2] ;
   wire \regIn[0][1] ;
   wire \regIn[0][0] ;
   wire \regIn[1][15] ;
   wire \regIn[1][14] ;
   wire \regIn[1][13] ;
   wire \regIn[1][12] ;
   wire \regIn[1][11] ;
   wire \regIn[1][10] ;
   wire \regIn[1][9] ;
   wire \regIn[1][8] ;
   wire \regIn[1][7] ;
   wire \regIn[1][6] ;
   wire \regIn[1][5] ;
   wire \regIn[1][4] ;
   wire \regIn[1][3] ;
   wire \regIn[1][2] ;
   wire \regIn[1][1] ;
   wire \regIn[1][0] ;
   wire \regIn[2][15] ;
   wire \regIn[2][14] ;
   wire \regIn[2][13] ;
   wire \regIn[2][12] ;
   wire \regIn[2][11] ;
   wire \regIn[2][10] ;
   wire \regIn[2][9] ;
   wire \regIn[2][8] ;
   wire \regIn[2][7] ;
   wire \regIn[2][6] ;
   wire \regIn[2][5] ;
   wire \regIn[2][4] ;
   wire \regIn[2][3] ;
   wire \regIn[2][2] ;
   wire \regIn[2][1] ;
   wire \regIn[2][0] ;
   wire \regIn[3][15] ;
   wire \regIn[3][14] ;
   wire \regIn[3][13] ;
   wire \regIn[3][12] ;
   wire \regIn[3][11] ;
   wire \regIn[3][10] ;
   wire \regIn[3][9] ;
   wire \regIn[3][8] ;
   wire \regIn[3][7] ;
   wire \regIn[3][6] ;
   wire \regIn[3][5] ;
   wire \regIn[3][4] ;
   wire \regIn[3][3] ;
   wire \regIn[3][2] ;
   wire \regIn[3][1] ;
   wire \regIn[3][0] ;
   wire \regIn[4][15] ;
   wire \regIn[4][14] ;
   wire \regIn[4][13] ;
   wire \regIn[4][12] ;
   wire \regIn[4][11] ;
   wire \regIn[4][10] ;
   wire \regIn[4][9] ;
   wire \regIn[4][8] ;
   wire \regIn[4][7] ;
   wire \regIn[4][6] ;
   wire \regIn[4][5] ;
   wire \regIn[4][4] ;
   wire \regIn[4][3] ;
   wire \regIn[4][2] ;
   wire \regIn[4][1] ;
   wire \regIn[4][0] ;
   wire \regIn[5][15] ;
   wire \regIn[5][14] ;
   wire \regIn[5][13] ;
   wire \regIn[5][12] ;
   wire \regIn[5][11] ;
   wire \regIn[5][10] ;
   wire \regIn[5][9] ;
   wire \regIn[5][8] ;
   wire \regIn[5][7] ;
   wire \regIn[5][6] ;
   wire \regIn[5][5] ;
   wire \regIn[5][4] ;
   wire \regIn[5][3] ;
   wire \regIn[5][2] ;
   wire \regIn[5][1] ;
   wire \regIn[5][0] ;
   wire \regIn[6][15] ;
   wire \regIn[6][14] ;
   wire \regIn[6][13] ;
   wire \regIn[6][12] ;
   wire \regIn[6][11] ;
   wire \regIn[6][10] ;
   wire \regIn[6][9] ;
   wire \regIn[6][8] ;
   wire \regIn[6][7] ;
   wire \regIn[6][6] ;
   wire \regIn[6][5] ;
   wire \regIn[6][4] ;
   wire \regIn[6][3] ;
   wire \regIn[6][2] ;
   wire \regIn[6][1] ;
   wire \regIn[6][0] ;
   wire \regIn[7][15] ;
   wire \regIn[7][14] ;
   wire \regIn[7][13] ;
   wire \regIn[7][12] ;
   wire \regIn[7][11] ;
   wire \regIn[7][10] ;
   wire \regIn[7][9] ;
   wire \regIn[7][8] ;
   wire \regIn[7][7] ;
   wire \regIn[7][6] ;
   wire \regIn[7][5] ;
   wire \regIn[7][4] ;
   wire \regIn[7][3] ;
   wire \regIn[7][2] ;
   wire \regIn[7][1] ;
   wire \regIn[7][0] ;
   wire \regIn[8][15] ;
   wire \regIn[8][14] ;
   wire \regIn[8][13] ;
   wire \regIn[8][12] ;
   wire \regIn[8][11] ;
   wire \regIn[8][10] ;
   wire \regIn[8][9] ;
   wire \regIn[8][8] ;
   wire \regIn[8][7] ;
   wire \regIn[8][6] ;
   wire \regIn[8][5] ;
   wire \regIn[8][4] ;
   wire \regIn[8][3] ;
   wire \regIn[8][2] ;
   wire \regIn[8][1] ;
   wire \regIn[8][0] ;
   wire \regIn[9][15] ;
   wire \regIn[9][14] ;
   wire \regIn[9][13] ;
   wire \regIn[9][12] ;
   wire \regIn[9][11] ;
   wire \regIn[9][10] ;
   wire \regIn[9][9] ;
   wire \regIn[9][8] ;
   wire \regIn[9][7] ;
   wire \regIn[9][6] ;
   wire \regIn[9][5] ;
   wire \regIn[9][4] ;
   wire \regIn[9][3] ;
   wire \regIn[9][2] ;
   wire \regIn[9][1] ;
   wire \regIn[9][0] ;
   wire \regIn[10][15] ;
   wire \regIn[10][14] ;
   wire \regIn[10][13] ;
   wire \regIn[10][12] ;
   wire \regIn[10][11] ;
   wire \regIn[10][10] ;
   wire \regIn[10][9] ;
   wire \regIn[10][8] ;
   wire \regIn[10][7] ;
   wire \regIn[10][6] ;
   wire \regIn[10][5] ;
   wire \regIn[10][4] ;
   wire \regIn[10][3] ;
   wire \regIn[10][2] ;
   wire \regIn[10][1] ;
   wire \regIn[10][0] ;
   wire \regIn[11][15] ;
   wire \regIn[11][14] ;
   wire \regIn[11][13] ;
   wire \regIn[11][12] ;
   wire \regIn[11][11] ;
   wire \regIn[11][10] ;
   wire \regIn[11][9] ;
   wire \regIn[11][8] ;
   wire \regIn[11][7] ;
   wire \regIn[11][6] ;
   wire \regIn[11][5] ;
   wire \regIn[11][4] ;
   wire \regIn[11][3] ;
   wire \regIn[11][2] ;
   wire \regIn[11][1] ;
   wire \regIn[11][0] ;
   wire \regIn[12][15] ;
   wire \regIn[12][14] ;
   wire \regIn[12][13] ;
   wire \regIn[12][12] ;
   wire \regIn[12][11] ;
   wire \regIn[12][10] ;
   wire \regIn[12][9] ;
   wire \regIn[12][8] ;
   wire \regIn[12][7] ;
   wire \regIn[12][6] ;
   wire \regIn[12][5] ;
   wire \regIn[12][4] ;
   wire \regIn[12][3] ;
   wire \regIn[12][2] ;
   wire \regIn[12][1] ;
   wire \regIn[12][0] ;
   wire \regIn[13][15] ;
   wire \regIn[13][14] ;
   wire \regIn[13][13] ;
   wire \regIn[13][12] ;
   wire \regIn[13][11] ;
   wire \regIn[13][10] ;
   wire \regIn[13][9] ;
   wire \regIn[13][8] ;
   wire \regIn[13][7] ;
   wire \regIn[13][6] ;
   wire \regIn[13][5] ;
   wire \regIn[13][4] ;
   wire \regIn[13][3] ;
   wire \regIn[13][2] ;
   wire \regIn[13][1] ;
   wire \regIn[13][0] ;
   wire \regIn[14][15] ;
   wire \regIn[14][14] ;
   wire \regIn[14][13] ;
   wire \regIn[14][12] ;
   wire \regIn[14][11] ;
   wire \regIn[14][10] ;
   wire \regIn[14][9] ;
   wire \regIn[14][8] ;
   wire \regIn[14][7] ;
   wire \regIn[14][6] ;
   wire \regIn[14][5] ;
   wire \regIn[14][4] ;
   wire \regIn[14][3] ;
   wire \regIn[14][2] ;
   wire \regIn[14][1] ;
   wire \regIn[14][0] ;
   wire \regIn[15][15] ;
   wire \regIn[15][14] ;
   wire \regIn[15][13] ;
   wire \regIn[15][12] ;
   wire \regIn[15][11] ;
   wire \regIn[15][10] ;
   wire \regIn[15][9] ;
   wire \regIn[15][8] ;
   wire \regIn[15][7] ;
   wire \regIn[15][6] ;
   wire \regIn[15][5] ;
   wire \regIn[15][4] ;
   wire \regIn[15][3] ;
   wire \regIn[15][2] ;
   wire \regIn[15][1] ;
   wire \regIn[15][0] ;
   wire \regIn[16][15] ;
   wire \regIn[16][14] ;
   wire \regIn[16][13] ;
   wire \regIn[16][12] ;
   wire \regIn[16][11] ;
   wire \regIn[16][10] ;
   wire \regIn[16][9] ;
   wire \regIn[16][8] ;
   wire \regIn[16][7] ;
   wire \regIn[16][6] ;
   wire \regIn[16][5] ;
   wire \regIn[16][4] ;
   wire \regIn[16][3] ;
   wire \regIn[16][2] ;
   wire \regIn[16][1] ;
   wire \regIn[16][0] ;
   wire \regIn[17][15] ;
   wire \regIn[17][14] ;
   wire \regIn[17][13] ;
   wire \regIn[17][12] ;
   wire \regIn[17][11] ;
   wire \regIn[17][10] ;
   wire \regIn[17][9] ;
   wire \regIn[17][8] ;
   wire \regIn[17][7] ;
   wire \regIn[17][6] ;
   wire \regIn[17][5] ;
   wire \regIn[17][4] ;
   wire \regIn[17][3] ;
   wire \regIn[17][2] ;
   wire \regIn[17][1] ;
   wire \regIn[17][0] ;
   wire \regIn[18][15] ;
   wire \regIn[18][14] ;
   wire \regIn[18][13] ;
   wire \regIn[18][12] ;
   wire \regIn[18][11] ;
   wire \regIn[18][10] ;
   wire \regIn[18][9] ;
   wire \regIn[18][8] ;
   wire \regIn[18][7] ;
   wire \regIn[18][6] ;
   wire \regIn[18][5] ;
   wire \regIn[18][4] ;
   wire \regIn[18][3] ;
   wire \regIn[18][2] ;
   wire \regIn[18][1] ;
   wire \regIn[18][0] ;
   wire \regIn[19][15] ;
   wire \regIn[19][14] ;
   wire \regIn[19][13] ;
   wire \regIn[19][12] ;
   wire \regIn[19][11] ;
   wire \regIn[19][10] ;
   wire \regIn[19][9] ;
   wire \regIn[19][8] ;
   wire \regIn[19][7] ;
   wire \regIn[19][6] ;
   wire \regIn[19][5] ;
   wire \regIn[19][4] ;
   wire \regIn[19][3] ;
   wire \regIn[19][2] ;
   wire \regIn[19][1] ;
   wire \regIn[19][0] ;
   wire \regIn[20][15] ;
   wire \regIn[20][14] ;
   wire \regIn[20][13] ;
   wire \regIn[20][12] ;
   wire \regIn[20][11] ;
   wire \regIn[20][10] ;
   wire \regIn[20][9] ;
   wire \regIn[20][8] ;
   wire \regIn[20][7] ;
   wire \regIn[20][6] ;
   wire \regIn[20][5] ;
   wire \regIn[20][4] ;
   wire \regIn[20][3] ;
   wire \regIn[20][2] ;
   wire \regIn[20][1] ;
   wire \regIn[20][0] ;
   wire \regIn[21][15] ;
   wire \regIn[21][14] ;
   wire \regIn[21][13] ;
   wire \regIn[21][12] ;
   wire \regIn[21][11] ;
   wire \regIn[21][10] ;
   wire \regIn[21][9] ;
   wire \regIn[21][8] ;
   wire \regIn[21][7] ;
   wire \regIn[21][6] ;
   wire \regIn[21][5] ;
   wire \regIn[21][4] ;
   wire \regIn[21][3] ;
   wire \regIn[21][2] ;
   wire \regIn[21][1] ;
   wire \regIn[21][0] ;
   wire \regIn[22][15] ;
   wire \regIn[22][14] ;
   wire \regIn[22][13] ;
   wire \regIn[22][12] ;
   wire \regIn[22][11] ;
   wire \regIn[22][10] ;
   wire \regIn[22][9] ;
   wire \regIn[22][8] ;
   wire \regIn[22][7] ;
   wire \regIn[22][6] ;
   wire \regIn[22][5] ;
   wire \regIn[22][4] ;
   wire \regIn[22][3] ;
   wire \regIn[22][2] ;
   wire \regIn[22][1] ;
   wire \regIn[22][0] ;
   wire \regIn[23][15] ;
   wire \regIn[23][14] ;
   wire \regIn[23][13] ;
   wire \regIn[23][12] ;
   wire \regIn[23][11] ;
   wire \regIn[23][10] ;
   wire \regIn[23][9] ;
   wire \regIn[23][8] ;
   wire \regIn[23][7] ;
   wire \regIn[23][6] ;
   wire \regIn[23][5] ;
   wire \regIn[23][4] ;
   wire \regIn[23][3] ;
   wire \regIn[23][2] ;
   wire \regIn[23][1] ;
   wire \regIn[23][0] ;
   wire \regIn[24][15] ;
   wire \regIn[24][14] ;
   wire \regIn[24][13] ;
   wire \regIn[24][12] ;
   wire \regIn[24][11] ;
   wire \regIn[24][10] ;
   wire \regIn[24][9] ;
   wire \regIn[24][8] ;
   wire \regIn[24][7] ;
   wire \regIn[24][6] ;
   wire \regIn[24][5] ;
   wire \regIn[24][4] ;
   wire \regIn[24][3] ;
   wire \regIn[24][2] ;
   wire \regIn[24][1] ;
   wire \regIn[24][0] ;
   wire \regIn[25][15] ;
   wire \regIn[25][14] ;
   wire \regIn[25][13] ;
   wire \regIn[25][12] ;
   wire \regIn[25][11] ;
   wire \regIn[25][10] ;
   wire \regIn[25][9] ;
   wire \regIn[25][8] ;
   wire \regIn[25][7] ;
   wire \regIn[25][6] ;
   wire \regIn[25][5] ;
   wire \regIn[25][4] ;
   wire \regIn[25][3] ;
   wire \regIn[25][2] ;
   wire \regIn[25][1] ;
   wire \regIn[25][0] ;
   wire \regIn[26][15] ;
   wire \regIn[26][14] ;
   wire \regIn[26][13] ;
   wire \regIn[26][12] ;
   wire \regIn[26][11] ;
   wire \regIn[26][10] ;
   wire \regIn[26][9] ;
   wire \regIn[26][8] ;
   wire \regIn[26][7] ;
   wire \regIn[26][6] ;
   wire \regIn[26][5] ;
   wire \regIn[26][4] ;
   wire \regIn[26][3] ;
   wire \regIn[26][2] ;
   wire \regIn[26][1] ;
   wire \regIn[26][0] ;
   wire \regIn[27][15] ;
   wire \regIn[27][14] ;
   wire \regIn[27][13] ;
   wire \regIn[27][12] ;
   wire \regIn[27][11] ;
   wire \regIn[27][10] ;
   wire \regIn[27][9] ;
   wire \regIn[27][8] ;
   wire \regIn[27][7] ;
   wire \regIn[27][6] ;
   wire \regIn[27][5] ;
   wire \regIn[27][4] ;
   wire \regIn[27][3] ;
   wire \regIn[27][2] ;
   wire \regIn[27][1] ;
   wire \regIn[27][0] ;
   wire \regIn[28][15] ;
   wire \regIn[28][14] ;
   wire \regIn[28][13] ;
   wire \regIn[28][12] ;
   wire \regIn[28][11] ;
   wire \regIn[28][10] ;
   wire \regIn[28][9] ;
   wire \regIn[28][8] ;
   wire \regIn[28][7] ;
   wire \regIn[28][6] ;
   wire \regIn[28][5] ;
   wire \regIn[28][4] ;
   wire \regIn[28][3] ;
   wire \regIn[28][2] ;
   wire \regIn[28][1] ;
   wire \regIn[28][0] ;
   wire \regIn[29][15] ;
   wire \regIn[29][14] ;
   wire \regIn[29][13] ;
   wire \regIn[29][12] ;
   wire \regIn[29][11] ;
   wire \regIn[29][10] ;
   wire \regIn[29][9] ;
   wire \regIn[29][8] ;
   wire \regIn[29][7] ;
   wire \regIn[29][6] ;
   wire \regIn[29][5] ;
   wire \regIn[29][4] ;
   wire \regIn[29][3] ;
   wire \regIn[29][2] ;
   wire \regIn[29][1] ;
   wire \regIn[29][0] ;
   wire \regIn[30][15] ;
   wire \regIn[30][14] ;
   wire \regIn[30][13] ;
   wire \regIn[30][12] ;
   wire \regIn[30][11] ;
   wire \regIn[30][10] ;
   wire \regIn[30][9] ;
   wire \regIn[30][8] ;
   wire \regIn[30][7] ;
   wire \regIn[30][6] ;
   wire \regIn[30][5] ;
   wire \regIn[30][4] ;
   wire \regIn[30][3] ;
   wire \regIn[30][2] ;
   wire \regIn[30][1] ;
   wire \regIn[30][0] ;
   wire \regIn[31][15] ;
   wire \regIn[31][14] ;
   wire \regIn[31][13] ;
   wire \regIn[31][12] ;
   wire \regIn[31][11] ;
   wire \regIn[31][10] ;
   wire \regIn[31][9] ;
   wire \regIn[31][8] ;
   wire \regIn[31][7] ;
   wire \regIn[31][6] ;
   wire \regIn[31][5] ;
   wire \regIn[31][4] ;
   wire \regIn[31][3] ;
   wire \regIn[31][2] ;
   wire \regIn[31][1] ;
   wire \regIn[31][0] ;
   wire N195;
   wire N196;
   wire N197;
   wire N198;
   wire N199;
   wire N200;
   wire N202;
   wire N203;
   wire N204;
   wire N205;
   wire N206;
   wire N207;
   wire N208;
   wire N209;
   wire N210;
   wire N211;
   wire N212;
   wire N213;
   wire N215;
   wire N216;
   wire N217;
   wire N218;
   wire N219;
   wire N220;
   wire N222;
   wire N223;
   wire N224;
   wire N225;
   wire N226;
   wire N228;
   wire N229;
   wire N230;
   wire N231;
   wire N232;
   wire N234;
   wire N235;
   wire N236;
   wire N237;
   wire N238;
   wire N240;
   wire N241;
   wire N242;
   wire N243;
   wire N244;
   wire N245;
   wire N247;
   wire N248;
   wire N249;
   wire N250;
   wire N251;
   wire N253;
   wire N254;
   wire N255;
   wire N256;
   wire N257;
   wire N259;
   wire N260;
   wire N261;
   wire N262;
   wire N263;
   wire N265;
   wire N266;
   wire N267;
   wire N268;
   wire N269;
   wire N271;
   wire N272;
   wire N273;
   wire N274;
   wire N275;
   wire N277;
   wire N278;
   wire N279;
   wire N280;
   wire N281;
   wire N283;
   wire N284;
   wire N285;
   wire N286;
   wire N287;
   wire N289;
   wire N290;
   wire N291;
   wire N292;
   wire N293;
   wire N296;
   wire N297;
   wire N298;
   wire N299;
   wire N300;
   wire N302;
   wire N303;
   wire N304;
   wire N305;
   wire N306;
   wire N307;
   wire N308;
   wire N309;
   wire N310;
   wire N311;
   wire N312;
   wire N314;
   wire N315;
   wire N316;
   wire N317;
   wire N318;
   wire N320;
   wire N321;
   wire N322;
   wire N323;
   wire N324;
   wire N326;
   wire N327;
   wire N328;
   wire N329;
   wire N330;
   wire N332;
   wire N333;
   wire N334;
   wire N335;
   wire N336;
   wire N338;
   wire N339;
   wire N340;
   wire N341;
   wire N342;
   wire N345;
   wire N346;
   wire N347;
   wire N348;
   wire N351;
   wire N352;
   wire N353;
   wire N354;
   wire N357;
   wire N358;
   wire N359;
   wire N360;
   wire N363;
   wire N364;
   wire N365;
   wire N366;
   wire N370;
   wire N371;
   wire N372;
   wire N376;
   wire N377;
   wire N378;
   wire N383;
   wire N384;
   wire N386;
   wire N387;
   wire N388;
   wire N389;
   wire N390;
   wire n2;
   wire n3;
   wire n4;
   wire n5;
   wire n6;
   wire n7;
   wire n8;
   wire n9;
   wire n10;
   wire n11;
   wire n12;
   wire n13;
   wire n14;
   wire n15;
   wire n16;
   wire n17;
   wire n18;
   wire n19;
   wire n20;
   wire n21;
   wire n22;
   wire n23;
   wire n24;
   wire n25;
   wire n26;
   wire n27;
   wire n28;
   wire n29;
   wire n30;
   wire n31;
   wire n32;
   wire n33;
   wire n34;
   wire n35;
   wire n36;
   wire n37;
   wire n38;
   wire n39;
   wire n40;
   wire n41;
   wire n42;
   wire n43;
   wire n44;
   wire n45;
   wire n46;
   wire n47;
   wire n48;
   wire n49;
   wire n50;
   wire n51;
   wire n52;
   wire n53;
   wire n54;
   wire n55;
   wire n56;
   wire n57;
   wire n58;
   wire n59;
   wire n60;
   wire n61;
   wire n62;
   wire n63;
   wire n64;
   wire n65;
   wire n66;
   wire n67;
   wire n68;
   wire n69;
   wire n70;
   wire n71;
   wire n72;
   wire n73;
   wire n74;
   wire n75;
   wire n76;
   wire n77;
   wire n78;
   wire n79;
   wire n80;
   wire n81;
   wire n82;
   wire n83;
   wire n84;
   wire n85;
   wire n86;
   wire n87;
   wire n88;
   wire n89;
   wire n90;
   wire n91;
   wire n92;
   wire n93;
   wire n94;
   wire n95;
   wire n96;
   wire n97;
   wire n98;
   wire n99;
   wire n100;
   wire n101;
   wire n102;
   wire n103;
   wire n104;
   wire n105;
   wire n106;
   wire n107;
   wire n108;
   wire n109;
   wire n110;
   wire n111;
   wire n112;
   wire n113;
   wire n114;
   wire n115;
   wire n116;
   wire n117;
   wire n118;
   wire n119;
   wire n120;
   wire n121;
   wire n122;
   wire n123;
   wire n124;
   wire n125;
   wire n126;
   wire n127;
   wire n128;
   wire n129;
   wire n130;
   wire n131;
   wire n132;
   wire n133;
   wire n134;
   wire n135;
   wire n136;
   wire n137;
   wire n138;
   wire n139;
   wire n140;
   wire n141;
   wire n142;
   wire n143;
   wire n144;
   wire n145;
   wire n146;
   wire n147;
   wire n148;
   wire n149;
   wire n150;
   wire n151;
   wire n152;
   wire n153;
   wire n154;
   wire n155;
   wire n156;
   wire n157;
   wire n158;
   wire n159;
   wire n160;
   wire n161;
   wire n162;
   wire n163;
   wire n164;
   wire n165;
   wire n166;
   wire n167;
   wire n168;
   wire n169;
   wire n170;
   wire n171;
   wire n172;
   wire n173;
   wire n174;
   wire n175;
   wire n176;
   wire n177;
   wire n178;
   wire n179;
   wire n180;
   wire n181;
   wire n182;
   wire n183;
   wire n184;
   wire n185;
   wire n186;
   wire n187;
   wire n188;
   wire n189;
   wire n190;
   wire n191;
   wire n192;
   wire n193;
   wire n194;
   wire n195;
   wire n196;
   wire n197;
   wire n198;
   wire n199;
   wire n200;
   wire n201;
   wire n202;
   wire n203;
   wire n204;
   wire n205;
   wire n206;
   wire n207;
   wire n208;
   wire n209;
   wire n210;
   wire n211;
   wire n212;
   wire n213;
   wire n214;
   wire n215;
   wire n216;
   wire n217;
   wire n218;
   wire n219;
   wire n220;
   wire n221;
   wire n222;
   wire n223;
   wire n224;
   wire n225;
   wire n226;
   wire n227;
   wire n228;
   wire n229;
   wire n230;
   wire n231;
   wire n232;
   wire n233;
   wire n234;
   wire n235;
   wire n236;
   wire n237;
   wire n238;
   wire n239;
   wire n240;
   wire n241;
   wire n242;
   wire n243;
   wire n244;
   wire n245;
   wire n246;
   wire n247;
   wire n248;
   wire n249;
   wire n250;
   wire n251;
   wire n252;
   wire n253;
   wire n254;
   wire n255;
   wire n256;
   wire n257;
   wire n258;
   wire n259;
   wire n260;
   wire n261;
   wire n262;
   wire n263;
   wire n264;
   wire n265;
   wire n266;
   wire n267;
   wire n268;
   wire n269;
   wire n270;
   wire n271;
   wire n272;
   wire n273;
   wire n274;
   wire n275;
   wire n276;
   wire n277;
   wire n278;
   wire n279;
   wire n280;
   wire n281;
   wire n282;
   wire n283;
   wire n284;
   wire n285;
   wire n286;
   wire n287;
   wire n288;
   wire n289;
   wire n290;
   wire n291;
   wire n292;
   wire n293;
   wire n294;
   wire n295;
   wire n296;
   wire n297;
   wire n298;
   wire n299;
   wire n300;
   wire n301;
   wire n302;
   wire n303;
   wire n304;
   wire n305;
   wire n306;
   wire n307;
   wire n308;
   wire n309;
   wire n310;
   wire n311;
   wire n312;
   wire n313;
   wire n314;
   wire n315;
   wire n316;
   wire n317;
   wire n318;
   wire n319;
   wire n320;
   wire n321;
   wire n322;
   wire n323;
   wire n324;
   wire n325;
   wire n326;
   wire n327;
   wire n328;
   wire n329;
   wire n330;
   wire n331;
   wire n332;
   wire n333;
   wire n334;
   wire n335;
   wire n336;
   wire n337;
   wire n338;
   wire n339;
   wire n340;
   wire n341;
   wire n342;
   wire n343;
   wire n344;
   wire n345;
   wire n346;
   wire n347;
   wire n348;
   wire n349;
   wire n350;
   wire n351;
   wire n352;
   wire n353;
   wire n354;
   wire n355;
   wire n356;
   wire n357;
   wire n358;
   wire n359;
   wire n360;
   wire n361;
   wire n362;
   wire n363;
   wire n364;
   wire n365;
   wire n366;
   wire n367;
   wire n368;
   wire n369;
   wire n370;
   wire n371;
   wire n372;
   wire n373;
   wire n374;
   wire n375;
   wire n376;
   wire n377;
   wire n378;
   wire n379;
   wire n380;
   wire n381;
   wire n382;
   wire n383;
   wire n384;
   wire n385;
   wire n386;
   wire n387;
   wire n388;
   wire n389;
   wire n390;
   wire n391;
   wire n392;
   wire n393;
   wire n394;
   wire n395;
   wire n396;
   wire n397;
   wire n398;
   wire n399;
   wire n400;
   wire n401;
   wire n402;
   wire n403;
   wire n404;
   wire n405;
   wire n406;
   wire n407;
   wire n408;
   wire n409;
   wire n410;
   wire n411;
   wire n412;
   wire n413;
   wire n414;
   wire n415;
   wire n416;
   wire n417;
   wire n418;
   wire n419;
   wire n420;
   wire n421;
   wire n422;
   wire n423;
   wire n424;
   wire n425;
   wire n426;
   wire n427;
   wire n428;
   wire n429;
   wire n430;
   wire n431;
   wire n432;
   wire n433;
   wire n434;
   wire n435;
   wire n436;
   wire n437;
   wire n438;
   wire n439;
   wire n440;
   wire n441;
   wire n442;
   wire n443;
   wire n444;
   wire n445;
   wire n446;
   wire n447;
   wire n448;
   wire n449;
   wire n450;
   wire n451;
   wire n452;
   wire n453;
   wire n454;
   wire n455;
   wire n456;
   wire n457;
   wire n458;
   wire n459;
   wire n460;
   wire n461;
   wire n462;
   wire n463;
   wire n464;
   wire n465;
   wire n466;
   wire n467;
   wire n468;
   wire n469;
   wire n470;
   wire n471;
   wire n472;
   wire n473;
   wire n474;
   wire n475;
   wire n476;
   wire n477;
   wire n478;
   wire n479;
   wire n480;
   wire n481;
   wire n482;
   wire n483;
   wire n484;
   wire n485;
   wire n486;
   wire n487;
   wire n488;
   wire n489;
   wire n490;
   wire n491;
   wire n492;
   wire n493;
   wire n494;
   wire n495;
   wire n496;
   wire n497;
   wire n498;
   wire n499;
   wire n500;
   wire n501;
   wire n502;
   wire n503;
   wire n504;
   wire n505;
   wire n506;
   wire n507;
   wire n508;
   wire n509;
   wire n510;
   wire n511;
   wire n512;
   wire n513;
   wire n514;
   wire n515;
   wire n516;
   wire n517;
   wire n518;
   wire n519;
   wire n520;
   wire n521;
   wire n522;
   wire n523;
   wire n524;
   wire n525;
   wire n526;
   wire n527;
   wire n528;
   wire n529;
   wire n530;
   wire n531;
   wire n532;
   wire n533;
   wire n534;
   wire n535;
   wire n536;
   wire n537;
   wire n538;
   wire n539;
   wire n540;
   wire n541;
   wire n542;
   wire n543;
   wire n544;
   wire n545;
   wire n546;
   wire n547;
   wire n548;
   wire n549;
   wire n550;
   wire n551;
   wire n552;
   wire n553;
   wire n554;
   wire n555;
   wire n556;
   wire n557;
   wire n558;
   wire n559;
   wire n560;
   wire n561;
   wire n562;
   wire n563;
   wire n564;
   wire n565;
   wire n566;
   wire n567;
   wire n568;
   wire n569;
   wire n570;
   wire n571;
   wire n572;
   wire n573;
   wire n574;
   wire n575;
   wire n576;
   wire n577;
   wire n578;
   wire n579;
   wire n580;
   wire n581;
   wire n582;
   wire n583;
   wire n584;
   wire n585;
   wire n586;
   wire n587;
   wire n588;
   wire n589;
   wire n590;
   wire n591;
   wire n592;
   wire n593;
   wire n594;
   wire n595;
   wire n596;
   wire n597;
   wire n598;
   wire n599;
   wire n600;
   wire n601;
   wire n602;
   wire n603;
   wire n604;
   wire n605;
   wire n606;
   wire n607;
   wire n608;
   wire n609;
   wire n610;
   wire n611;
   wire n612;
   wire n613;
   wire n614;
   wire n615;
   wire n616;
   wire n617;
   wire n618;
   wire n619;
   wire n620;
   wire n621;
   wire n622;
   wire n623;
   wire n624;
   wire n625;
   wire n626;
   wire n627;
   wire n628;
   wire n629;
   wire n630;
   wire n631;
   wire n632;
   wire n633;
   wire n634;
   wire n635;
   wire n636;
   wire n637;
   wire n638;
   wire n639;
   wire n640;
   wire n641;
   wire n642;
   wire n643;
   wire n644;
   wire n645;
   wire n646;
   wire n647;
   wire n648;
   wire n649;
   wire n650;
   wire n651;
   wire n652;
   wire n653;
   wire n654;
   wire n655;
   wire n656;
   wire n657;
   wire n658;
   wire n659;
   wire n660;
   wire n661;
   wire n662;
   wire n663;
   wire n664;
   wire n665;
   wire n666;
   wire n667;
   wire n668;
   wire n669;
   wire n670;
   wire n671;
   wire n672;
   wire n673;
   wire n674;
   wire n675;
   wire n676;
   wire n677;
   wire n678;
   wire n679;
   wire n680;
   wire n681;
   wire n682;
   wire n683;
   wire n684;
   wire n685;
   wire n686;
   wire n687;
   wire n688;
   wire n689;
   wire n690;
   wire n691;
   wire n692;
   wire n693;
   wire n694;
   wire n695;
   wire n696;
   wire n697;
   wire n698;
   wire n699;
   wire n700;
   wire n701;
   wire n702;
   wire n703;
   wire n704;
   wire n705;
   wire n706;
   wire n707;
   wire n708;
   wire n709;
   wire n710;
   wire n711;
   wire n712;
   wire n713;
   wire n714;
   wire n715;
   wire n716;
   wire n717;
   wire n718;
   wire n719;
   wire n720;
   wire n721;
   wire n722;
   wire n723;
   wire n724;
   wire n725;
   wire n726;
   wire n727;
   wire n728;
   wire n729;
   wire n730;
   wire n731;
   wire n732;
   wire n733;
   wire n734;
   wire n735;
   wire n736;
   wire n737;
   wire n738;
   wire n739;
   wire n740;
   wire n741;
   wire n742;
   wire n743;
   wire n744;
   wire n745;
   wire n746;
   wire n747;
   wire n748;
   wire n749;
   wire n750;
   wire n751;
   wire n752;
   wire n753;
   wire n754;
   wire n755;
   wire n756;
   wire n757;
   wire n758;
   wire n759;
   wire n760;
   wire n761;
   wire n762;
   wire n763;
   wire n764;
   wire n765;
   wire n766;
   wire n767;
   wire n768;
   wire n769;
   wire n770;
   wire n771;
   wire n772;
   wire n773;
   wire n774;
   wire n775;
   wire n776;
   wire n777;
   wire n778;
   wire n779;
   wire n780;
   wire n781;
   wire n782;
   wire n783;
   wire n784;
   wire n785;
   wire n786;
   wire n787;
   wire n788;
   wire n789;
   wire n790;
   wire n791;
   wire n792;
   wire n793;
   wire n794;
   wire n795;
   wire n796;
   wire n797;
   wire n798;
   wire n799;
   wire n800;
   wire n801;
   wire n802;
   wire n803;
   wire n804;
   wire n805;
   wire n806;
   wire n807;
   wire n808;
   wire n809;
   wire n810;
   wire n811;
   wire n812;
   wire n813;
   wire n814;
   wire n815;
   wire n816;
   wire n817;
   wire n818;
   wire n819;
   wire n820;
   wire n821;
   wire n822;
   wire n823;
   wire n824;
   wire n825;
   wire n826;
   wire n827;
   wire n828;
   wire n829;
   wire n830;
   wire n831;
   wire n832;
   wire n833;
   wire n834;
   wire n835;
   wire n836;
   wire n837;
   wire n838;
   wire n839;
   wire n840;
   wire n841;
   wire n842;
   wire n843;
   wire n844;
   wire n845;
   wire n846;
   wire n847;
   wire n848;
   wire n849;
   wire n850;
   wire n851;
   wire n852;
   wire n853;
   wire n854;
   wire n855;
   wire n856;
   wire n857;
   wire n858;
   wire n859;
   wire n860;
   wire n861;
   wire n862;
   wire n863;
   wire n864;
   wire n865;
   wire n866;
   wire n867;
   wire n868;
   wire n869;
   wire n870;
   wire n871;
   wire n872;
   wire n873;
   wire n874;
   wire n875;
   wire n876;
   wire n877;
   wire n878;
   wire n879;
   wire n880;
   wire n881;
   wire n882;
   wire n883;
   wire n884;
   wire n885;
   wire n886;
   wire n887;
   wire n888;
   wire n889;
   wire n890;
   wire n891;
   wire n892;
   wire n893;
   wire n894;
   wire n895;
   wire n896;
   wire n897;
   wire n898;
   wire n899;
   wire n900;
   wire n901;
   wire n902;
   wire n903;
   wire n904;
   wire n905;
   wire n906;
   wire n907;
   wire n908;
   wire n909;
   wire n910;
   wire n911;
   wire n912;
   wire n913;
   wire n914;
   wire n915;
   wire n916;
   wire n917;
   wire n918;
   wire n919;
   wire n920;
   wire n921;
   wire n922;
   wire n923;
   wire n924;
   wire n925;
   wire n926;
   wire n927;
   wire n928;
   wire n929;
   wire n930;
   wire n931;
   wire n932;
   wire n933;
   wire n934;
   wire n935;
   wire n936;
   wire n937;
   wire n938;
   wire n939;
   wire n940;
   wire n941;
   wire n942;
   wire n943;
   wire n944;
   wire n945;
   wire n946;
   wire n947;
   wire n948;
   wire n949;
   wire n950;
   wire n951;
   wire n952;
   wire n953;
   wire n954;
   wire n955;
   wire n956;
   wire n957;
   wire n958;
   wire n959;
   wire n960;
   wire n961;
   wire n962;
   wire n963;
   wire n964;
   wire n965;
   wire n966;
   wire n967;
   wire n968;
   wire n969;
   wire n970;
   wire n971;
   wire n972;
   wire n973;
   wire n974;
   wire n975;
   wire n976;
   wire n977;
   wire n978;
   wire n979;
   wire n980;
   wire n981;
   wire n982;
   wire n983;
   wire n984;
   wire n985;
   wire n986;
   wire n987;
   wire n988;
   wire n989;
   wire n990;
   wire n991;
   wire n992;
   wire n993;
   wire n994;
   wire n995;
   wire n996;
   wire n997;
   wire n998;
   wire n999;
   wire n1000;
   wire n1001;
   wire n1002;
   wire n1003;
   wire n1004;
   wire n1005;
   wire n1006;
   wire n1007;
   wire n1008;
   wire n1009;
   wire n1010;
   wire n1011;
   wire n1012;
   wire n1013;
   wire n1014;
   wire n1015;
   wire n1016;
   wire n1017;
   wire n1018;
   wire n1019;
   wire n1020;
   wire n1021;
   wire n1022;
   wire n1023;
   wire n1024;
   wire n1025;
   wire n1026;
   wire n1027;
   wire n1028;
   wire n1029;
   wire n1030;
   wire n1031;
   wire n1032;
   wire n1033;
   wire n1034;
   wire n1035;
   wire n1036;
   wire n1037;
   wire n1038;
   wire n1039;
   wire n1040;
   wire n1041;
   wire n1042;
   wire n1043;
   wire n1044;
   wire n1045;
   wire n1046;
   wire n1047;
   wire n1048;
   wire n1049;
   wire n1050;
   wire n1051;
   wire n1052;
   wire n1053;
   wire n1054;
   wire n1055;
   wire n1056;
   wire n1057;
   wire n1058;
   wire n1059;
   wire n1060;
   wire n1061;
   wire n1062;
   wire n1063;
   wire n1064;
   wire n1065;
   wire n1066;
   wire n1067;
   wire n1068;
   wire n1069;
   wire n1070;
   wire n1071;
   wire n1072;
   wire n1073;
   wire n1074;
   wire n1075;
   wire n1076;
   wire n1077;
   wire n1078;
   wire n1079;
   wire n1080;
   wire n1081;
   wire n1082;
   wire n1083;
   wire n1084;
   wire n1085;
   wire n1086;
   wire n1087;
   wire n1088;
   wire n1089;
   wire n1090;
   wire n1091;
   wire n1092;
   wire n1093;
   wire n1094;
   wire n1095;
   wire n1096;
   wire n1097;
   wire n1098;
   wire n1099;
   wire n1100;
   wire n1101;
   wire n1102;
   wire n1103;
   wire n1104;
   wire n1105;
   wire n1106;
   wire n1107;
   wire n1108;
   wire n1109;
   wire n1110;
   wire n1111;
   wire n1112;
   wire n1113;
   wire n1114;
   wire n1115;
   wire n1116;
   wire n1117;
   wire n1118;
   wire n1119;
   wire n1120;
   wire n1121;
   wire n1122;
   wire n1123;
   wire n1124;
   wire n1125;
   wire n1126;
   wire n1127;
   wire n1128;
   wire n1129;
   wire n1130;
   wire n1131;
   wire n1132;
   wire n1133;
   wire n1134;
   wire n1135;
   wire n1136;
   wire n1137;
   wire n1138;
   wire n1139;
   wire n1140;
   wire n1141;
   wire n1142;
   wire n1143;
   wire n1144;
   wire n1145;
   wire n1146;
   wire n1147;
   wire n1148;
   wire n1149;
   wire n1150;
   wire n1151;
   wire n1152;
   wire n1153;
   wire n1154;
   wire n1155;
   wire n1156;
   wire n1157;
   wire n1158;
   wire n1159;
   wire n1160;
   wire n1161;
   wire n1162;
   wire n1163;
   wire n1164;
   wire n1165;
   wire n1166;
   wire n1167;
   wire n1168;
   wire n1169;
   wire n1170;
   wire n1171;
   wire n1172;
   wire n1173;
   wire n1174;
   wire n1175;
   wire n1176;
   wire n1177;
   wire n1178;
   wire n1179;
   wire n1180;
   wire n1181;
   wire n1182;
   wire n1183;
   wire n1184;
   wire n1185;
   wire n1186;
   wire n1187;
   wire n1188;
   wire n1189;
   wire n1190;
   wire n1191;
   wire n1192;
   wire n1193;
   wire n1194;
   wire n1195;
   wire n1196;
   wire n1197;
   wire n1198;
   wire n1199;
   wire n1200;
   wire n1201;
   wire n1202;
   wire n1203;
   wire n1204;
   wire n1205;
   wire n1206;
   wire n1207;
   wire n1208;
   wire n1209;
   wire n1210;
   wire n1211;
   wire n1212;
   wire n1213;
   wire n1214;
   wire n1215;
   wire n1216;
   wire n1217;
   wire n1218;
   wire n1219;
   wire n1220;
   wire n1221;
   wire n1222;
   wire n1223;
   wire n1224;
   wire n1225;
   wire n1226;
   wire n1227;
   wire n1228;
   wire n1229;
   wire n1230;
   wire n1231;
   wire n1232;
   wire n1233;
   wire n1234;
   wire n1235;
   wire n1236;
   wire n1237;
   wire n1238;
   wire n1239;
   wire n1240;
   wire n1241;
   wire n1271;

   assign N208 = addressIn[4] ;

   // Module instantiations
   CLKBUF_X3 clk__L2_I13 (
	.Z(clk__L2_N13),
	.A(clk__L1_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUF_X3 clk__L2_I12 (
	.Z(clk__L2_N12),
	.A(clk__L1_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUF_X3 clk__L2_I11 (
	.Z(clk__L2_N11),
	.A(clk__L1_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUF_X3 clk__L2_I10 (
	.Z(clk__L2_N10),
	.A(clk__L1_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUF_X3 clk__L2_I9 (
	.Z(clk__L2_N9),
	.A(clk__L1_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUF_X3 clk__L2_I8 (
	.Z(clk__L2_N8),
	.A(clk__L1_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUF_X3 clk__L2_I7 (
	.Z(clk__L2_N7),
	.A(clk__L1_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUF_X3 clk__L2_I6 (
	.Z(clk__L2_N6),
	.A(clk__L1_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUF_X3 clk__L2_I5 (
	.Z(clk__L2_N5),
	.A(clk__L1_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUF_X3 clk__L2_I4 (
	.Z(clk__L2_N4),
	.A(clk__L1_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUF_X3 clk__L2_I3 (
	.Z(clk__L2_N3),
	.A(clk__L1_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUF_X3 clk__L2_I2 (
	.Z(clk__L2_N2),
	.A(clk__L1_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUF_X3 clk__L2_I1 (
	.Z(clk__L2_N1),
	.A(clk__L1_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUF_X3 clk__L2_I0 (
	.Z(clk__L2_N0),
	.A(clk__L1_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUF_X3 clk__L1_I0 (
	.Z(clk__L1_N0),
	.A(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   BUF_X1 FE_OFC75_n569 (
	.Z(FE_OFN75_n569),
	.A(n569), 
	.VDD(VDD), 
	.VSS(VSS));
   BUF_X2 FE_OFC74_n568 (
	.Z(FE_OFN74_n568),
	.A(n568), 
	.VDD(VDD), 
	.VSS(VSS));
   BUF_X1 FE_OFC73_n574 (
	.Z(FE_OFN73_n574),
	.A(n574), 
	.VDD(VDD), 
	.VSS(VSS));
   BUF_X2 FE_OFC72_n573 (
	.Z(FE_OFN72_n573),
	.A(n573), 
	.VDD(VDD), 
	.VSS(VSS));
   BUF_X1 FE_OFC71_n603 (
	.Z(FE_OFN71_n603),
	.A(n603), 
	.VDD(VDD), 
	.VSS(VSS));
   BUF_X1 FE_OFC70_n602 (
	.Z(FE_OFN70_n602),
	.A(n602), 
	.VDD(VDD), 
	.VSS(VSS));
   BUF_X1 FE_OFC69_n608 (
	.Z(FE_OFN69_n608),
	.A(n608), 
	.VDD(VDD), 
	.VSS(VSS));
   BUF_X1 FE_OFC68_n607 (
	.Z(FE_OFN68_n607),
	.A(n607), 
	.VDD(VDD), 
	.VSS(VSS));
   BUF_X1 FE_OFC67_n579 (
	.Z(FE_OFN67_n579),
	.A(n579), 
	.VDD(VDD), 
	.VSS(VSS));
   BUF_X2 FE_OFC66_n578 (
	.Z(FE_OFN66_n578),
	.A(n578), 
	.VDD(VDD), 
	.VSS(VSS));
   BUF_X1 FE_OFC65_n584 (
	.Z(FE_OFN65_n584),
	.A(n584), 
	.VDD(VDD), 
	.VSS(VSS));
   BUF_X1 FE_OFC64_n583 (
	.Z(FE_OFN64_n583),
	.A(n583), 
	.VDD(VDD), 
	.VSS(VSS));
   BUF_X1 FE_OFC63_n593 (
	.Z(FE_OFN63_n593),
	.A(n593), 
	.VDD(VDD), 
	.VSS(VSS));
   BUF_X1 FE_OFC62_n592 (
	.Z(FE_OFN62_n592),
	.A(n592), 
	.VDD(VDD), 
	.VSS(VSS));
   BUF_X1 FE_OFC61_n598 (
	.Z(FE_OFN61_n598),
	.A(n598), 
	.VDD(VDD), 
	.VSS(VSS));
   BUF_X1 FE_OFC60_n597 (
	.Z(FE_OFN60_n597),
	.A(n597), 
	.VDD(VDD), 
	.VSS(VSS));
   BUF_X2 FE_OFC59_write (
	.Z(FE_OFN59_write),
	.A(FE_OFN40_write), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUF_X3 FE_OFC58_write (
	.Z(FE_OFN58_write),
	.A(FE_OFN40_write), 
	.VDD(VDD), 
	.VSS(VSS));
   BUF_X1 FE_OFC57_write (
	.Z(FE_OFN57_write),
	.A(FE_OFN40_write), 
	.VDD(VDD), 
	.VSS(VSS));
   BUF_X2 FE_OFC56_write (
	.Z(FE_OFN56_write),
	.A(FE_OFN40_write), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUF_X3 FE_OFC55_write (
	.Z(FE_OFN55_write),
	.A(FE_OFN38_write), 
	.VDD(VDD), 
	.VSS(VSS));
   BUF_X1 FE_OFC54_write (
	.Z(FE_OFN54_write),
	.A(FE_OFN40_write), 
	.VDD(VDD), 
	.VSS(VSS));
   BUF_X1 FE_OFC53_write (
	.Z(FE_OFN53_write),
	.A(FE_OFN40_write), 
	.VDD(VDD), 
	.VSS(VSS));
   BUF_X1 FE_OFC51_write (
	.Z(FE_OFN51_write),
	.A(FE_OFN40_write), 
	.VDD(VDD), 
	.VSS(VSS));
   BUF_X1 FE_OFC50_write (
	.Z(FE_OFN50_write),
	.A(FE_OFN38_write), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUF_X2 FE_OFC49_write (
	.Z(FE_OFN49_write),
	.A(FE_OFN40_write), 
	.VDD(VDD), 
	.VSS(VSS));
   BUF_X1 FE_OFC48_write (
	.Z(FE_OFN48_write),
	.A(FE_OFN26_write), 
	.VDD(VDD), 
	.VSS(VSS));
   BUF_X1 FE_OFC47_write (
	.Z(FE_OFN47_write),
	.A(FE_OFN40_write), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUF_X3 FE_OFC46_write (
	.Z(FE_OFN46_write),
	.A(FE_OFN26_write), 
	.VDD(VDD), 
	.VSS(VSS));
   BUF_X1 FE_OFC45_write (
	.Z(FE_OFN45_write),
	.A(FE_OFN38_write), 
	.VDD(VDD), 
	.VSS(VSS));
   BUF_X4 FE_OFC44_write (
	.Z(FE_OFN44_write),
	.A(FE_OFN32_write), 
	.VDD(VDD), 
	.VSS(VSS));
   BUF_X1 FE_OFC43_write (
	.Z(FE_OFN43_write),
	.A(FE_OFN40_write), 
	.VDD(VDD), 
	.VSS(VSS));
   BUF_X1 FE_OFC42_write (
	.Z(FE_OFN42_write),
	.A(FE_OFN26_write), 
	.VDD(VDD), 
	.VSS(VSS));
   BUF_X2 FE_OFC41_write (
	.Z(FE_OFN41_write),
	.A(FE_OFN32_write), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUF_X3 FE_OFC40_write (
	.Z(FE_OFN40_write),
	.A(FE_OFN21_write), 
	.VDD(VDD), 
	.VSS(VSS));
   BUF_X1 FE_OFC39_write (
	.Z(FE_OFN39_write),
	.A(FE_OFN26_write), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUF_X3 FE_OFC38_write (
	.Z(FE_OFN38_write),
	.A(FE_OFN21_write), 
	.VDD(VDD), 
	.VSS(VSS));
   BUF_X1 FE_OFC35_write (
	.Z(FE_OFN35_write),
	.A(FE_OFN26_write), 
	.VDD(VDD), 
	.VSS(VSS));
   BUF_X1 FE_OFC34_write (
	.Z(FE_OFN34_write),
	.A(FE_OFN21_write), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUF_X2 FE_OFC32_write (
	.Z(FE_OFN32_write),
	.A(FE_OFN21_write), 
	.VDD(VDD), 
	.VSS(VSS));
   BUF_X1 FE_OFC31_write (
	.Z(FE_OFN31_write),
	.A(FE_OFN21_write), 
	.VDD(VDD), 
	.VSS(VSS));
   BUF_X1 FE_OFC30_write (
	.Z(FE_OFN30_write),
	.A(FE_OFN26_write), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUF_X1 FE_OFC29_write (
	.Z(FE_OFN29_write),
	.A(FE_OFN21_write), 
	.VDD(VDD), 
	.VSS(VSS));
   BUF_X2 FE_OFC28_write (
	.Z(FE_OFN28_write),
	.A(FE_OFN26_write), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUF_X3 FE_OFC26_write (
	.Z(FE_OFN26_write),
	.A(FE_OFN18_write), 
	.VDD(VDD), 
	.VSS(VSS));
   BUF_X1 FE_OFC25_write (
	.Z(FE_OFN25_write),
	.A(FE_OFN21_write), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUF_X1 FE_OFC24_write (
	.Z(FE_OFN24_write),
	.A(FE_OFN21_write), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUF_X1 FE_OFC23_write (
	.Z(FE_OFN23_write),
	.A(FE_OFN18_write), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUF_X1 FE_OFC22_write (
	.Z(FE_OFN22_write),
	.A(FE_OFN21_write), 
	.VDD(VDD), 
	.VSS(VSS));
   BUF_X32 FE_OFC21_write (
	.Z(FE_OFN21_write),
	.A(write), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUF_X1 FE_OFC20_write (
	.Z(FE_OFN20_write),
	.A(write), 
	.VDD(VDD), 
	.VSS(VSS));
   BUF_X16 FE_OFC18_write (
	.Z(FE_OFN18_write),
	.A(write), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUF_X1 FE_OFC17_write (
	.Z(FE_OFN17_write),
	.A(write), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUF_X2 FE_OFC16_write (
	.Z(FE_OFN16_write),
	.A(FE_OFN15_write), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUF_X1 FE_OFC15_write (
	.Z(FE_OFN15_write),
	.A(write), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 I_36 (
	.ZN(N390),
	.A(N389), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2_X1 C1077 (
	.ZN(N389),
	.A2(N388),
	.A1(N200), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2_X1 C1076 (
	.ZN(N388),
	.A2(N387),
	.A1(N207), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2_X1 C1075 (
	.ZN(N387),
	.A2(N386),
	.A1(N220), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2_X1 C1074 (
	.ZN(N386),
	.A2(N307),
	.A1(N245), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 I_35 (
	.ZN(N384),
	.A(N383), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 I_34 (
	.ZN(N378),
	.A(N377), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2_X1 C1056 (
	.ZN(N377),
	.A2(N376),
	.A1(N200), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 I_33 (
	.ZN(N372),
	.A(N371), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 I_32 (
	.ZN(N366),
	.A(N365), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2_X1 C1037 (
	.ZN(N365),
	.A2(N364),
	.A1(N200), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2_X1 C1036 (
	.ZN(N364),
	.A2(N363),
	.A1(N207), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 I_31 (
	.ZN(N360),
	.A(N359), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2_X1 C1026 (
	.ZN(N358),
	.A2(N357),
	.A1(N207), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 I_30 (
	.ZN(N354),
	.A(N353), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2_X1 C1018 (
	.ZN(N353),
	.A2(N352),
	.A1(N200), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 I_29 (
	.ZN(N348),
	.A(N347), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 I_28 (
	.ZN(N342),
	.A(N341), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2_X1 C1001 (
	.ZN(N341),
	.A2(N340),
	.A1(N200), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2_X1 C1000 (
	.ZN(N340),
	.A2(N339),
	.A1(N207), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2_X1 C999 (
	.ZN(N339),
	.A2(N338),
	.A1(N220), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 I_27 (
	.ZN(N336),
	.A(N335), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2_X1 C990 (
	.ZN(N334),
	.A2(N333),
	.A1(N207), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2_X1 C989 (
	.ZN(N333),
	.A2(N332),
	.A1(N220), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 I_26 (
	.ZN(N330),
	.A(N329), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2_X1 C982 (
	.ZN(N329),
	.A2(N328),
	.A1(N200), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2_X1 C980 (
	.ZN(N327),
	.A2(N326),
	.A1(N220), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 I_25 (
	.ZN(N324),
	.A(N323), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2_X1 C971 (
	.ZN(N321),
	.A2(N320),
	.A1(N220), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 I_24 (
	.ZN(N318),
	.A(N317), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2_X1 C965 (
	.ZN(N317),
	.A2(N316),
	.A1(N200), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2_X1 C964 (
	.ZN(N316),
	.A2(N315),
	.A1(N207), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 I_23 (
	.ZN(N312),
	.A(N311), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2_X1 C955 (
	.ZN(N310),
	.A2(N309),
	.A1(N207), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 I_22 (
	.ZN(N306),
	.A(N305), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2_X1 C948 (
	.ZN(N305),
	.A2(N304),
	.A1(N200), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 I_21 (
	.ZN(N300),
	.A(N299), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 I_20 (
	.ZN(N307),
	.A(n1271), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 I_19 (
	.ZN(N293),
	.A(N292), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2_X1 C933 (
	.ZN(N292),
	.A2(N291),
	.A1(N200), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2_X1 C932 (
	.ZN(N291),
	.A2(N290),
	.A1(N207), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2_X1 C931 (
	.ZN(N290),
	.A2(N289),
	.A1(N220), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 I_18 (
	.ZN(N287),
	.A(N286), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2_X1 C922 (
	.ZN(N285),
	.A2(N284),
	.A1(N207), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2_X1 C921 (
	.ZN(N284),
	.A2(N283),
	.A1(N220), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 I_17 (
	.ZN(N281),
	.A(N280), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2_X1 C914 (
	.ZN(N280),
	.A2(N279),
	.A1(N200), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2_X1 C912 (
	.ZN(N278),
	.A2(N277),
	.A1(N220), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 I_16 (
	.ZN(N275),
	.A(N274), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2_X1 C903 (
	.ZN(N272),
	.A2(N271),
	.A1(N220), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 I_15 (
	.ZN(N269),
	.A(N268), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2_X1 C897 (
	.ZN(N268),
	.A2(N267),
	.A1(N200), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2_X1 C896 (
	.ZN(N267),
	.A2(N266),
	.A1(N207), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 I_14 (
	.ZN(N263),
	.A(N262), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2_X1 C887 (
	.ZN(N261),
	.A2(N260),
	.A1(N207), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 I_13 (
	.ZN(N257),
	.A(N256), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2_X1 C880 (
	.ZN(N256),
	.A2(N255),
	.A1(N200), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 I_12 (
	.ZN(N251),
	.A(N250), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 I_10 (
	.ZN(N244),
	.A(N243), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2_X1 C865 (
	.ZN(N243),
	.A2(N242),
	.A1(N200), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2_X1 C864 (
	.ZN(N242),
	.A2(N241),
	.A1(N207), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2_X1 C863 (
	.ZN(N241),
	.A2(N240),
	.A1(N220), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 I_9 (
	.ZN(N238),
	.A(N237), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2_X1 C855 (
	.ZN(N236),
	.A2(N235),
	.A1(N207), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2_X1 C854 (
	.ZN(N235),
	.A2(N234),
	.A1(N220), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 I_8 (
	.ZN(N232),
	.A(N231), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2_X1 C848 (
	.ZN(N231),
	.A2(N230),
	.A1(N200), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2_X1 C846 (
	.ZN(N229),
	.A2(N228),
	.A1(N220), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 I_7 (
	.ZN(N226),
	.A(N225), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2_X1 C838 (
	.ZN(N223),
	.A2(N222),
	.A1(N220), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 I_5 (
	.ZN(N219),
	.A(N218), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2_X1 C833 (
	.ZN(N218),
	.A2(N217),
	.A1(N200), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2_X1 C832 (
	.ZN(N217),
	.A2(N216),
	.A1(N207), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 I_4 (
	.ZN(N213),
	.A(N212), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2_X1 C824 (
	.ZN(N211),
	.A2(N210),
	.A1(N207), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 I_2 (
	.ZN(N206),
	.A(N205), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2_X1 C818 (
	.ZN(N205),
	.A2(N204),
	.A1(N200), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 I_0 (
	.ZN(N199),
	.A(N198), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U2 (
	.ZN(\regIn[9][9] ),
	.B2(n4),
	.B1(N257),
	.A2(n3),
	.A1(n2), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U3 (
	.ZN(\regIn[9][8] ),
	.B2(n6),
	.B1(N257),
	.A2(n5),
	.A1(n2), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U4 (
	.ZN(\regIn[9][7] ),
	.B2(n8),
	.B1(N257),
	.A2(n7),
	.A1(n2), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U5 (
	.ZN(\regIn[9][6] ),
	.B2(n10),
	.B1(N257),
	.A2(n9),
	.A1(n2), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U6 (
	.ZN(\regIn[9][5] ),
	.B2(n12),
	.B1(N257),
	.A2(n11),
	.A1(n2), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U7 (
	.ZN(\regIn[9][4] ),
	.B2(n14),
	.B1(N257),
	.A2(n13),
	.A1(n2), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U8 (
	.ZN(\regIn[9][3] ),
	.B2(n16),
	.B1(N257),
	.A2(n15),
	.A1(n2), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U9 (
	.ZN(\regIn[9][2] ),
	.B2(n18),
	.B1(N257),
	.A2(n17),
	.A1(n2), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U10 (
	.ZN(\regIn[9][1] ),
	.B2(n20),
	.B1(N257),
	.A2(n19),
	.A1(n2), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U11 (
	.ZN(\regIn[9][15] ),
	.B2(n22),
	.B1(N257),
	.A2(n21),
	.A1(n2), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U12 (
	.ZN(\regIn[9][14] ),
	.B2(n24),
	.B1(N257),
	.A2(n23),
	.A1(n2), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U13 (
	.ZN(\regIn[9][13] ),
	.B2(n26),
	.B1(N257),
	.A2(n25),
	.A1(n2), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U14 (
	.ZN(\regIn[9][12] ),
	.B2(n28),
	.B1(N257),
	.A2(n27),
	.A1(n2), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U15 (
	.ZN(\regIn[9][11] ),
	.B2(n30),
	.B1(N257),
	.A2(n29),
	.A1(n2), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U16 (
	.ZN(\regIn[9][10] ),
	.B2(n32),
	.B1(N257),
	.A2(n31),
	.A1(n2), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U17 (
	.ZN(\regIn[9][0] ),
	.B2(n34),
	.B1(N257),
	.A2(n33),
	.A1(n2), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U18 (
	.ZN(n2),
	.A(N257), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U19 (
	.ZN(\regIn[8][9] ),
	.B2(n36),
	.B1(N251),
	.A2(n35),
	.A1(n3), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U20 (
	.ZN(\regIn[8][8] ),
	.B2(n37),
	.B1(N251),
	.A2(n35),
	.A1(n5), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U21 (
	.ZN(\regIn[8][7] ),
	.B2(n38),
	.B1(N251),
	.A2(n35),
	.A1(n7), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U22 (
	.ZN(\regIn[8][6] ),
	.B2(n39),
	.B1(N251),
	.A2(n35),
	.A1(n9), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U23 (
	.ZN(\regIn[8][5] ),
	.B2(n40),
	.B1(N251),
	.A2(n35),
	.A1(n11), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U24 (
	.ZN(\regIn[8][4] ),
	.B2(n41),
	.B1(N251),
	.A2(n35),
	.A1(n13), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U25 (
	.ZN(\regIn[8][3] ),
	.B2(n42),
	.B1(N251),
	.A2(n35),
	.A1(n15), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U26 (
	.ZN(\regIn[8][2] ),
	.B2(n43),
	.B1(N251),
	.A2(n35),
	.A1(n17), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U27 (
	.ZN(\regIn[8][1] ),
	.B2(n44),
	.B1(N251),
	.A2(n35),
	.A1(n19), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U28 (
	.ZN(\regIn[8][15] ),
	.B2(n45),
	.B1(N251),
	.A2(n35),
	.A1(n21), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U29 (
	.ZN(\regIn[8][14] ),
	.B2(n46),
	.B1(N251),
	.A2(n35),
	.A1(n23), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U30 (
	.ZN(\regIn[8][13] ),
	.B2(n47),
	.B1(N251),
	.A2(n35),
	.A1(n25), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U31 (
	.ZN(\regIn[8][12] ),
	.B2(n48),
	.B1(N251),
	.A2(n35),
	.A1(n27), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U32 (
	.ZN(\regIn[8][11] ),
	.B2(n49),
	.B1(N251),
	.A2(n35),
	.A1(n29), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U33 (
	.ZN(\regIn[8][10] ),
	.B2(n50),
	.B1(N251),
	.A2(n35),
	.A1(n31), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U34 (
	.ZN(\regIn[8][0] ),
	.B2(n51),
	.B1(N251),
	.A2(n35),
	.A1(n33), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U35 (
	.ZN(n35),
	.A(N251), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U36 (
	.ZN(\regIn[7][9] ),
	.A(n52), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U37 (
	.ZN(n52),
	.B2(\regOut[7][9] ),
	.B1(n53),
	.A2(N244),
	.A1(dataIn[9]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U38 (
	.ZN(\regIn[7][8] ),
	.A(n54), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U39 (
	.ZN(n54),
	.B2(\regOut[7][8] ),
	.B1(n53),
	.A2(N244),
	.A1(dataIn[8]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U40 (
	.ZN(\regIn[7][7] ),
	.A(n55), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U41 (
	.ZN(n55),
	.B2(\regOut[7][7] ),
	.B1(n53),
	.A2(N244),
	.A1(dataIn[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U42 (
	.ZN(\regIn[7][6] ),
	.A(n56), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U43 (
	.ZN(n56),
	.B2(\regOut[7][6] ),
	.B1(n53),
	.A2(N244),
	.A1(dataIn[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U44 (
	.ZN(\regIn[7][5] ),
	.A(n57), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U45 (
	.ZN(n57),
	.B2(\regOut[7][5] ),
	.B1(n53),
	.A2(N244),
	.A1(dataIn[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U46 (
	.ZN(\regIn[7][4] ),
	.A(n58), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U47 (
	.ZN(n58),
	.B2(\regOut[7][4] ),
	.B1(n53),
	.A2(N244),
	.A1(dataIn[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U48 (
	.ZN(\regIn[7][3] ),
	.A(n59), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U49 (
	.ZN(n59),
	.B2(\regOut[7][3] ),
	.B1(n53),
	.A2(N244),
	.A1(dataIn[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U50 (
	.ZN(\regIn[7][2] ),
	.A(n60), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U51 (
	.ZN(n60),
	.B2(\regOut[7][2] ),
	.B1(n53),
	.A2(N244),
	.A1(dataIn[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U52 (
	.ZN(\regIn[7][1] ),
	.A(n61), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U53 (
	.ZN(n61),
	.B2(\regOut[7][1] ),
	.B1(n53),
	.A2(N244),
	.A1(dataIn[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U54 (
	.ZN(\regIn[7][15] ),
	.A(n62), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U55 (
	.ZN(n62),
	.B2(\regOut[7][15] ),
	.B1(n53),
	.A2(N244),
	.A1(dataIn[15]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U56 (
	.ZN(\regIn[7][14] ),
	.A(n63), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U57 (
	.ZN(n63),
	.B2(\regOut[7][14] ),
	.B1(n53),
	.A2(N244),
	.A1(dataIn[14]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U58 (
	.ZN(\regIn[7][13] ),
	.A(n64), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U59 (
	.ZN(n64),
	.B2(\regOut[7][13] ),
	.B1(n53),
	.A2(N244),
	.A1(dataIn[13]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U60 (
	.ZN(\regIn[7][12] ),
	.A(n65), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U61 (
	.ZN(n65),
	.B2(\regOut[7][12] ),
	.B1(n53),
	.A2(N244),
	.A1(dataIn[12]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U62 (
	.ZN(\regIn[7][11] ),
	.A(n66), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U63 (
	.ZN(n66),
	.B2(\regOut[7][11] ),
	.B1(n53),
	.A2(N244),
	.A1(dataIn[11]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U64 (
	.ZN(\regIn[7][10] ),
	.A(n67), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U65 (
	.ZN(n67),
	.B2(\regOut[7][10] ),
	.B1(n53),
	.A2(N244),
	.A1(dataIn[10]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U66 (
	.ZN(\regIn[7][0] ),
	.A(n68), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U67 (
	.ZN(n68),
	.B2(\regOut[7][0] ),
	.B1(n53),
	.A2(N244),
	.A1(dataIn[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U68 (
	.ZN(n53),
	.A(N244), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U69 (
	.ZN(\regIn[6][9] ),
	.A(n69), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U70 (
	.ZN(n69),
	.B2(\regOut[6][9] ),
	.B1(n70),
	.A2(N238),
	.A1(dataIn[9]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U71 (
	.ZN(\regIn[6][8] ),
	.A(n71), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U72 (
	.ZN(n71),
	.B2(\regOut[6][8] ),
	.B1(n70),
	.A2(N238),
	.A1(dataIn[8]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U73 (
	.ZN(\regIn[6][7] ),
	.A(n72), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U74 (
	.ZN(n72),
	.B2(\regOut[6][7] ),
	.B1(n70),
	.A2(N238),
	.A1(dataIn[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U75 (
	.ZN(\regIn[6][6] ),
	.A(n73), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U76 (
	.ZN(n73),
	.B2(\regOut[6][6] ),
	.B1(n70),
	.A2(N238),
	.A1(dataIn[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U77 (
	.ZN(\regIn[6][5] ),
	.A(n74), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U78 (
	.ZN(n74),
	.B2(\regOut[6][5] ),
	.B1(n70),
	.A2(N238),
	.A1(dataIn[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U79 (
	.ZN(\regIn[6][4] ),
	.A(n75), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U80 (
	.ZN(n75),
	.B2(\regOut[6][4] ),
	.B1(n70),
	.A2(N238),
	.A1(dataIn[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U81 (
	.ZN(\regIn[6][3] ),
	.A(n76), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U82 (
	.ZN(n76),
	.B2(\regOut[6][3] ),
	.B1(n70),
	.A2(N238),
	.A1(dataIn[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U83 (
	.ZN(\regIn[6][2] ),
	.A(n77), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U84 (
	.ZN(n77),
	.B2(\regOut[6][2] ),
	.B1(n70),
	.A2(N238),
	.A1(dataIn[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U85 (
	.ZN(\regIn[6][1] ),
	.A(n78), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U86 (
	.ZN(n78),
	.B2(\regOut[6][1] ),
	.B1(n70),
	.A2(N238),
	.A1(dataIn[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U87 (
	.ZN(\regIn[6][15] ),
	.A(n79), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U88 (
	.ZN(n79),
	.B2(\regOut[6][15] ),
	.B1(n70),
	.A2(N238),
	.A1(dataIn[15]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U89 (
	.ZN(\regIn[6][14] ),
	.A(n80), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U90 (
	.ZN(n80),
	.B2(\regOut[6][14] ),
	.B1(n70),
	.A2(N238),
	.A1(dataIn[14]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U91 (
	.ZN(\regIn[6][13] ),
	.A(n81), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U92 (
	.ZN(n81),
	.B2(\regOut[6][13] ),
	.B1(n70),
	.A2(N238),
	.A1(dataIn[13]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U93 (
	.ZN(\regIn[6][12] ),
	.A(n82), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U94 (
	.ZN(n82),
	.B2(\regOut[6][12] ),
	.B1(n70),
	.A2(N238),
	.A1(dataIn[12]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U95 (
	.ZN(\regIn[6][11] ),
	.A(n83), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U96 (
	.ZN(n83),
	.B2(\regOut[6][11] ),
	.B1(n70),
	.A2(N238),
	.A1(dataIn[11]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U97 (
	.ZN(\regIn[6][10] ),
	.A(n84), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U98 (
	.ZN(n84),
	.B2(\regOut[6][10] ),
	.B1(n70),
	.A2(N238),
	.A1(dataIn[10]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U99 (
	.ZN(\regIn[6][0] ),
	.A(n85), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U100 (
	.ZN(n85),
	.B2(\regOut[6][0] ),
	.B1(n70),
	.A2(N238),
	.A1(dataIn[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U101 (
	.ZN(n70),
	.A(N238), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U102 (
	.ZN(\regIn[5][9] ),
	.B2(n87),
	.B1(N232),
	.A2(n86),
	.A1(n3), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U103 (
	.ZN(\regIn[5][8] ),
	.B2(n88),
	.B1(N232),
	.A2(n86),
	.A1(n5), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U104 (
	.ZN(\regIn[5][7] ),
	.B2(n89),
	.B1(N232),
	.A2(n86),
	.A1(n7), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U105 (
	.ZN(\regIn[5][6] ),
	.B2(n90),
	.B1(N232),
	.A2(n86),
	.A1(n9), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U106 (
	.ZN(\regIn[5][5] ),
	.B2(n91),
	.B1(N232),
	.A2(n86),
	.A1(n11), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U107 (
	.ZN(\regIn[5][4] ),
	.B2(n92),
	.B1(N232),
	.A2(n86),
	.A1(n13), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U108 (
	.ZN(\regIn[5][3] ),
	.B2(n93),
	.B1(N232),
	.A2(n86),
	.A1(n15), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U109 (
	.ZN(\regIn[5][2] ),
	.B2(n94),
	.B1(N232),
	.A2(n86),
	.A1(n17), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U110 (
	.ZN(\regIn[5][1] ),
	.B2(n95),
	.B1(N232),
	.A2(n86),
	.A1(n19), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U111 (
	.ZN(\regIn[5][15] ),
	.B2(n96),
	.B1(N232),
	.A2(n86),
	.A1(n21), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U112 (
	.ZN(\regIn[5][14] ),
	.B2(n97),
	.B1(N232),
	.A2(n86),
	.A1(n23), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U113 (
	.ZN(\regIn[5][13] ),
	.B2(n98),
	.B1(N232),
	.A2(n86),
	.A1(n25), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U114 (
	.ZN(\regIn[5][12] ),
	.B2(n99),
	.B1(N232),
	.A2(n86),
	.A1(n27), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U115 (
	.ZN(\regIn[5][11] ),
	.B2(n100),
	.B1(N232),
	.A2(n86),
	.A1(n29), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U116 (
	.ZN(\regIn[5][10] ),
	.B2(n101),
	.B1(N232),
	.A2(n86),
	.A1(n31), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U117 (
	.ZN(\regIn[5][0] ),
	.B2(n102),
	.B1(N232),
	.A2(n86),
	.A1(n33), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U118 (
	.ZN(n86),
	.A(N232), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U119 (
	.ZN(\regIn[4][9] ),
	.B2(n104),
	.B1(N226),
	.A2(n103),
	.A1(n3), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U120 (
	.ZN(\regIn[4][8] ),
	.B2(n105),
	.B1(N226),
	.A2(n103),
	.A1(n5), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U121 (
	.ZN(\regIn[4][7] ),
	.B2(n106),
	.B1(N226),
	.A2(n103),
	.A1(n7), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U122 (
	.ZN(\regIn[4][6] ),
	.B2(n107),
	.B1(N226),
	.A2(n103),
	.A1(n9), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U123 (
	.ZN(\regIn[4][5] ),
	.B2(n108),
	.B1(N226),
	.A2(n103),
	.A1(n11), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U124 (
	.ZN(\regIn[4][4] ),
	.B2(n109),
	.B1(N226),
	.A2(n103),
	.A1(n13), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U125 (
	.ZN(\regIn[4][3] ),
	.B2(n110),
	.B1(N226),
	.A2(n103),
	.A1(n15), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U126 (
	.ZN(\regIn[4][2] ),
	.B2(n111),
	.B1(N226),
	.A2(n103),
	.A1(n17), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U127 (
	.ZN(\regIn[4][1] ),
	.B2(n112),
	.B1(N226),
	.A2(n103),
	.A1(n19), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U128 (
	.ZN(\regIn[4][15] ),
	.B2(n113),
	.B1(N226),
	.A2(n103),
	.A1(n21), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U129 (
	.ZN(\regIn[4][14] ),
	.B2(n114),
	.B1(N226),
	.A2(n103),
	.A1(n23), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U130 (
	.ZN(\regIn[4][13] ),
	.B2(n115),
	.B1(N226),
	.A2(n103),
	.A1(n25), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U131 (
	.ZN(\regIn[4][12] ),
	.B2(n116),
	.B1(N226),
	.A2(n103),
	.A1(n27), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U132 (
	.ZN(\regIn[4][11] ),
	.B2(n117),
	.B1(N226),
	.A2(n103),
	.A1(n29), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U133 (
	.ZN(\regIn[4][10] ),
	.B2(n118),
	.B1(N226),
	.A2(n103),
	.A1(n31), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U134 (
	.ZN(\regIn[4][0] ),
	.B2(n119),
	.B1(N226),
	.A2(n103),
	.A1(n33), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U135 (
	.ZN(n103),
	.A(N226), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U136 (
	.ZN(\regIn[3][9] ),
	.A(n120), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U137 (
	.ZN(n120),
	.B2(\regOut[3][9] ),
	.B1(n121),
	.A2(N219),
	.A1(dataIn[9]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U138 (
	.ZN(\regIn[3][8] ),
	.A(n122), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U139 (
	.ZN(n122),
	.B2(\regOut[3][8] ),
	.B1(n121),
	.A2(N219),
	.A1(dataIn[8]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U140 (
	.ZN(\regIn[3][7] ),
	.A(n123), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U141 (
	.ZN(n123),
	.B2(\regOut[3][7] ),
	.B1(n121),
	.A2(N219),
	.A1(dataIn[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U142 (
	.ZN(\regIn[3][6] ),
	.A(n124), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U143 (
	.ZN(n124),
	.B2(\regOut[3][6] ),
	.B1(n121),
	.A2(N219),
	.A1(dataIn[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U144 (
	.ZN(\regIn[3][5] ),
	.A(n125), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U145 (
	.ZN(n125),
	.B2(\regOut[3][5] ),
	.B1(n121),
	.A2(N219),
	.A1(dataIn[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U146 (
	.ZN(\regIn[3][4] ),
	.A(n126), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U147 (
	.ZN(n126),
	.B2(\regOut[3][4] ),
	.B1(n121),
	.A2(N219),
	.A1(dataIn[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U148 (
	.ZN(\regIn[3][3] ),
	.A(n127), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U149 (
	.ZN(n127),
	.B2(\regOut[3][3] ),
	.B1(n121),
	.A2(N219),
	.A1(dataIn[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U150 (
	.ZN(\regIn[3][2] ),
	.A(n128), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U151 (
	.ZN(n128),
	.B2(\regOut[3][2] ),
	.B1(n121),
	.A2(N219),
	.A1(dataIn[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U152 (
	.ZN(\regIn[3][1] ),
	.A(n129), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U153 (
	.ZN(n129),
	.B2(\regOut[3][1] ),
	.B1(n121),
	.A2(N219),
	.A1(dataIn[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U154 (
	.ZN(\regIn[3][15] ),
	.A(n130), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U155 (
	.ZN(n130),
	.B2(\regOut[3][15] ),
	.B1(n121),
	.A2(N219),
	.A1(dataIn[15]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U156 (
	.ZN(\regIn[3][14] ),
	.A(n131), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U157 (
	.ZN(n131),
	.B2(\regOut[3][14] ),
	.B1(n121),
	.A2(N219),
	.A1(dataIn[14]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U158 (
	.ZN(\regIn[3][13] ),
	.A(n132), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U159 (
	.ZN(n132),
	.B2(\regOut[3][13] ),
	.B1(n121),
	.A2(N219),
	.A1(dataIn[13]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U160 (
	.ZN(\regIn[3][12] ),
	.A(n133), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U161 (
	.ZN(n133),
	.B2(\regOut[3][12] ),
	.B1(n121),
	.A2(N219),
	.A1(dataIn[12]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U162 (
	.ZN(\regIn[3][11] ),
	.A(n134), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U163 (
	.ZN(n134),
	.B2(\regOut[3][11] ),
	.B1(n121),
	.A2(N219),
	.A1(dataIn[11]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U164 (
	.ZN(\regIn[3][10] ),
	.A(n135), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U165 (
	.ZN(n135),
	.B2(\regOut[3][10] ),
	.B1(n121),
	.A2(N219),
	.A1(dataIn[10]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U166 (
	.ZN(\regIn[3][0] ),
	.A(n136), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U167 (
	.ZN(n136),
	.B2(\regOut[3][0] ),
	.B1(n121),
	.A2(N219),
	.A1(dataIn[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U168 (
	.ZN(n121),
	.A(N219), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U169 (
	.ZN(\regIn[31][9] ),
	.B2(n138),
	.B1(N390),
	.A2(n137),
	.A1(n3), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U170 (
	.ZN(\regIn[31][8] ),
	.B2(n139),
	.B1(N390),
	.A2(n137),
	.A1(n5), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U171 (
	.ZN(\regIn[31][7] ),
	.B2(n140),
	.B1(N390),
	.A2(n137),
	.A1(n7), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U172 (
	.ZN(\regIn[31][6] ),
	.B2(n141),
	.B1(N390),
	.A2(n137),
	.A1(n9), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U173 (
	.ZN(\regIn[31][5] ),
	.B2(n142),
	.B1(N390),
	.A2(n137),
	.A1(n11), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U174 (
	.ZN(\regIn[31][4] ),
	.B2(n143),
	.B1(N390),
	.A2(n137),
	.A1(n13), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U175 (
	.ZN(\regIn[31][3] ),
	.B2(n144),
	.B1(N390),
	.A2(n137),
	.A1(n15), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U176 (
	.ZN(\regIn[31][2] ),
	.B2(n145),
	.B1(N390),
	.A2(n137),
	.A1(n17), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U177 (
	.ZN(\regIn[31][1] ),
	.B2(n146),
	.B1(N390),
	.A2(n137),
	.A1(n19), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U178 (
	.ZN(\regIn[31][15] ),
	.B2(n147),
	.B1(N390),
	.A2(n137),
	.A1(n21), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U179 (
	.ZN(\regIn[31][14] ),
	.B2(n148),
	.B1(N390),
	.A2(n137),
	.A1(n23), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U180 (
	.ZN(\regIn[31][13] ),
	.B2(n149),
	.B1(N390),
	.A2(n137),
	.A1(n25), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U181 (
	.ZN(\regIn[31][12] ),
	.B2(n150),
	.B1(N390),
	.A2(n137),
	.A1(n27), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U182 (
	.ZN(\regIn[31][11] ),
	.B2(n151),
	.B1(N390),
	.A2(n137),
	.A1(n29), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U183 (
	.ZN(\regIn[31][10] ),
	.B2(n152),
	.B1(N390),
	.A2(n137),
	.A1(n31), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U184 (
	.ZN(\regIn[31][0] ),
	.B2(n153),
	.B1(N390),
	.A2(n137),
	.A1(n33), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U185 (
	.ZN(n137),
	.A(N390), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U186 (
	.ZN(\regIn[30][9] ),
	.B2(n155),
	.B1(N384),
	.A2(n154),
	.A1(n3), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U187 (
	.ZN(\regIn[30][8] ),
	.B2(n156),
	.B1(N384),
	.A2(n154),
	.A1(n5), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U188 (
	.ZN(\regIn[30][7] ),
	.B2(n157),
	.B1(N384),
	.A2(n154),
	.A1(n7), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U189 (
	.ZN(\regIn[30][6] ),
	.B2(n158),
	.B1(N384),
	.A2(n154),
	.A1(n9), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U190 (
	.ZN(\regIn[30][5] ),
	.B2(n159),
	.B1(N384),
	.A2(n154),
	.A1(n11), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U191 (
	.ZN(\regIn[30][4] ),
	.B2(n160),
	.B1(N384),
	.A2(n154),
	.A1(n13), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U192 (
	.ZN(\regIn[30][3] ),
	.B2(n161),
	.B1(N384),
	.A2(n154),
	.A1(n15), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U193 (
	.ZN(\regIn[30][2] ),
	.B2(n162),
	.B1(N384),
	.A2(n154),
	.A1(n17), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U194 (
	.ZN(\regIn[30][1] ),
	.B2(n163),
	.B1(N384),
	.A2(n154),
	.A1(n19), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U195 (
	.ZN(\regIn[30][15] ),
	.B2(n164),
	.B1(N384),
	.A2(n154),
	.A1(n21), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U196 (
	.ZN(\regIn[30][14] ),
	.B2(n165),
	.B1(N384),
	.A2(n154),
	.A1(n23), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U197 (
	.ZN(\regIn[30][13] ),
	.B2(n166),
	.B1(N384),
	.A2(n154),
	.A1(n25), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U198 (
	.ZN(\regIn[30][12] ),
	.B2(n167),
	.B1(N384),
	.A2(n154),
	.A1(n27), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U199 (
	.ZN(\regIn[30][11] ),
	.B2(n168),
	.B1(N384),
	.A2(n154),
	.A1(n29), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U200 (
	.ZN(\regIn[30][10] ),
	.B2(n169),
	.B1(N384),
	.A2(n154),
	.A1(n31), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U201 (
	.ZN(\regIn[30][0] ),
	.B2(n170),
	.B1(N384),
	.A2(n154),
	.A1(n33), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U202 (
	.ZN(n154),
	.A(N384), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U203 (
	.ZN(\regIn[2][9] ),
	.A(n171), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U204 (
	.ZN(n171),
	.B2(\regOut[2][9] ),
	.B1(n172),
	.A2(N213),
	.A1(dataIn[9]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U205 (
	.ZN(\regIn[2][8] ),
	.A(n173), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U206 (
	.ZN(n173),
	.B2(\regOut[2][8] ),
	.B1(n172),
	.A2(N213),
	.A1(dataIn[8]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U207 (
	.ZN(\regIn[2][7] ),
	.A(n174), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U208 (
	.ZN(n174),
	.B2(\regOut[2][7] ),
	.B1(n172),
	.A2(N213),
	.A1(dataIn[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U209 (
	.ZN(\regIn[2][6] ),
	.A(n175), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U210 (
	.ZN(n175),
	.B2(\regOut[2][6] ),
	.B1(n172),
	.A2(N213),
	.A1(dataIn[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U211 (
	.ZN(\regIn[2][5] ),
	.A(n176), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U212 (
	.ZN(n176),
	.B2(\regOut[2][5] ),
	.B1(n172),
	.A2(N213),
	.A1(dataIn[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U213 (
	.ZN(\regIn[2][4] ),
	.A(n177), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U214 (
	.ZN(n177),
	.B2(\regOut[2][4] ),
	.B1(n172),
	.A2(N213),
	.A1(dataIn[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U215 (
	.ZN(\regIn[2][3] ),
	.A(n178), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U216 (
	.ZN(n178),
	.B2(\regOut[2][3] ),
	.B1(n172),
	.A2(N213),
	.A1(dataIn[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U217 (
	.ZN(\regIn[2][2] ),
	.A(n179), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U218 (
	.ZN(n179),
	.B2(\regOut[2][2] ),
	.B1(n172),
	.A2(N213),
	.A1(dataIn[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U219 (
	.ZN(\regIn[2][1] ),
	.A(n180), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U220 (
	.ZN(n180),
	.B2(\regOut[2][1] ),
	.B1(n172),
	.A2(N213),
	.A1(dataIn[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U221 (
	.ZN(\regIn[2][15] ),
	.A(n181), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U222 (
	.ZN(n181),
	.B2(\regOut[2][15] ),
	.B1(n172),
	.A2(N213),
	.A1(dataIn[15]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U223 (
	.ZN(\regIn[2][14] ),
	.A(n182), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U224 (
	.ZN(n182),
	.B2(\regOut[2][14] ),
	.B1(n172),
	.A2(N213),
	.A1(dataIn[14]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U225 (
	.ZN(\regIn[2][13] ),
	.A(n183), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U226 (
	.ZN(n183),
	.B2(\regOut[2][13] ),
	.B1(n172),
	.A2(N213),
	.A1(dataIn[13]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U227 (
	.ZN(\regIn[2][12] ),
	.A(n184), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U228 (
	.ZN(n184),
	.B2(\regOut[2][12] ),
	.B1(n172),
	.A2(N213),
	.A1(dataIn[12]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U229 (
	.ZN(\regIn[2][11] ),
	.A(n185), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U230 (
	.ZN(n185),
	.B2(\regOut[2][11] ),
	.B1(n172),
	.A2(N213),
	.A1(dataIn[11]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U231 (
	.ZN(\regIn[2][10] ),
	.A(n186), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U232 (
	.ZN(n186),
	.B2(\regOut[2][10] ),
	.B1(n172),
	.A2(N213),
	.A1(dataIn[10]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U233 (
	.ZN(\regIn[2][0] ),
	.A(n187), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U234 (
	.ZN(n187),
	.B2(\regOut[2][0] ),
	.B1(n172),
	.A2(N213),
	.A1(dataIn[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U235 (
	.ZN(n172),
	.A(N213), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U236 (
	.ZN(\regIn[29][9] ),
	.A(n188), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U237 (
	.ZN(n188),
	.B2(\regOut[29][9] ),
	.B1(n189),
	.A2(N378),
	.A1(dataIn[9]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U238 (
	.ZN(\regIn[29][8] ),
	.A(n190), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U239 (
	.ZN(n190),
	.B2(\regOut[29][8] ),
	.B1(n189),
	.A2(N378),
	.A1(dataIn[8]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U240 (
	.ZN(\regIn[29][7] ),
	.A(n191), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U241 (
	.ZN(n191),
	.B2(\regOut[29][7] ),
	.B1(n189),
	.A2(N378),
	.A1(dataIn[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U242 (
	.ZN(\regIn[29][6] ),
	.A(n192), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U243 (
	.ZN(n192),
	.B2(\regOut[29][6] ),
	.B1(n189),
	.A2(N378),
	.A1(dataIn[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U244 (
	.ZN(\regIn[29][5] ),
	.A(n193), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U245 (
	.ZN(n193),
	.B2(\regOut[29][5] ),
	.B1(n189),
	.A2(N378),
	.A1(dataIn[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U246 (
	.ZN(\regIn[29][4] ),
	.A(n194), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U247 (
	.ZN(n194),
	.B2(\regOut[29][4] ),
	.B1(n189),
	.A2(N378),
	.A1(dataIn[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U248 (
	.ZN(\regIn[29][3] ),
	.A(n195), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U249 (
	.ZN(n195),
	.B2(\regOut[29][3] ),
	.B1(n189),
	.A2(N378),
	.A1(dataIn[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U250 (
	.ZN(\regIn[29][2] ),
	.A(n196), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U251 (
	.ZN(n196),
	.B2(\regOut[29][2] ),
	.B1(n189),
	.A2(N378),
	.A1(dataIn[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U252 (
	.ZN(\regIn[29][1] ),
	.A(n197), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U253 (
	.ZN(n197),
	.B2(\regOut[29][1] ),
	.B1(n189),
	.A2(N378),
	.A1(dataIn[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U254 (
	.ZN(\regIn[29][15] ),
	.A(n198), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U255 (
	.ZN(n198),
	.B2(\regOut[29][15] ),
	.B1(n189),
	.A2(N378),
	.A1(dataIn[15]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U256 (
	.ZN(\regIn[29][14] ),
	.A(n199), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U257 (
	.ZN(n199),
	.B2(\regOut[29][14] ),
	.B1(n189),
	.A2(N378),
	.A1(dataIn[14]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U258 (
	.ZN(\regIn[29][13] ),
	.A(n200), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U259 (
	.ZN(n200),
	.B2(\regOut[29][13] ),
	.B1(n189),
	.A2(N378),
	.A1(dataIn[13]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U260 (
	.ZN(\regIn[29][12] ),
	.A(n201), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U261 (
	.ZN(n201),
	.B2(\regOut[29][12] ),
	.B1(n189),
	.A2(N378),
	.A1(dataIn[12]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U262 (
	.ZN(\regIn[29][11] ),
	.A(n202), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U263 (
	.ZN(n202),
	.B2(\regOut[29][11] ),
	.B1(n189),
	.A2(N378),
	.A1(dataIn[11]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U264 (
	.ZN(\regIn[29][10] ),
	.A(n203), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U265 (
	.ZN(n203),
	.B2(\regOut[29][10] ),
	.B1(n189),
	.A2(N378),
	.A1(dataIn[10]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U266 (
	.ZN(\regIn[29][0] ),
	.A(n204), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U267 (
	.ZN(n204),
	.B2(\regOut[29][0] ),
	.B1(n189),
	.A2(N378),
	.A1(dataIn[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U268 (
	.ZN(n189),
	.A(N378), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U269 (
	.ZN(\regIn[28][9] ),
	.A(n205), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U270 (
	.ZN(n205),
	.B2(\regOut[28][9] ),
	.B1(n206),
	.A2(N372),
	.A1(dataIn[9]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U271 (
	.ZN(\regIn[28][8] ),
	.A(n207), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U272 (
	.ZN(n207),
	.B2(\regOut[28][8] ),
	.B1(n206),
	.A2(N372),
	.A1(dataIn[8]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U273 (
	.ZN(\regIn[28][7] ),
	.A(n208), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U274 (
	.ZN(n208),
	.B2(\regOut[28][7] ),
	.B1(n206),
	.A2(N372),
	.A1(dataIn[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U275 (
	.ZN(\regIn[28][6] ),
	.A(n209), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U276 (
	.ZN(n209),
	.B2(\regOut[28][6] ),
	.B1(n206),
	.A2(N372),
	.A1(dataIn[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U277 (
	.ZN(\regIn[28][5] ),
	.A(n210), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U278 (
	.ZN(n210),
	.B2(\regOut[28][5] ),
	.B1(n206),
	.A2(N372),
	.A1(dataIn[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U279 (
	.ZN(\regIn[28][4] ),
	.A(n211), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U280 (
	.ZN(n211),
	.B2(\regOut[28][4] ),
	.B1(n206),
	.A2(N372),
	.A1(dataIn[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U281 (
	.ZN(\regIn[28][3] ),
	.A(n212), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U282 (
	.ZN(n212),
	.B2(\regOut[28][3] ),
	.B1(n206),
	.A2(N372),
	.A1(dataIn[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U283 (
	.ZN(\regIn[28][2] ),
	.A(n213), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U284 (
	.ZN(n213),
	.B2(\regOut[28][2] ),
	.B1(n206),
	.A2(N372),
	.A1(dataIn[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U285 (
	.ZN(\regIn[28][1] ),
	.A(n214), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U286 (
	.ZN(n214),
	.B2(\regOut[28][1] ),
	.B1(n206),
	.A2(N372),
	.A1(dataIn[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U287 (
	.ZN(\regIn[28][15] ),
	.A(n215), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U288 (
	.ZN(n215),
	.B2(\regOut[28][15] ),
	.B1(n206),
	.A2(N372),
	.A1(dataIn[15]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U289 (
	.ZN(\regIn[28][14] ),
	.A(n216), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U290 (
	.ZN(n216),
	.B2(\regOut[28][14] ),
	.B1(n206),
	.A2(N372),
	.A1(dataIn[14]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U291 (
	.ZN(\regIn[28][13] ),
	.A(n217), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U292 (
	.ZN(n217),
	.B2(\regOut[28][13] ),
	.B1(n206),
	.A2(N372),
	.A1(dataIn[13]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U293 (
	.ZN(\regIn[28][12] ),
	.A(n218), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U294 (
	.ZN(n218),
	.B2(\regOut[28][12] ),
	.B1(n206),
	.A2(N372),
	.A1(dataIn[12]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U295 (
	.ZN(\regIn[28][11] ),
	.A(n219), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U296 (
	.ZN(n219),
	.B2(\regOut[28][11] ),
	.B1(n206),
	.A2(N372),
	.A1(dataIn[11]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U297 (
	.ZN(\regIn[28][10] ),
	.A(n220), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U298 (
	.ZN(n220),
	.B2(\regOut[28][10] ),
	.B1(n206),
	.A2(N372),
	.A1(dataIn[10]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U299 (
	.ZN(\regIn[28][0] ),
	.A(n221), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U300 (
	.ZN(n221),
	.B2(\regOut[28][0] ),
	.B1(n206),
	.A2(N372),
	.A1(dataIn[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U301 (
	.ZN(n206),
	.A(N372), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U302 (
	.ZN(\regIn[27][9] ),
	.A(n222), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U303 (
	.ZN(n222),
	.B2(\regOut[27][9] ),
	.B1(n223),
	.A2(N366),
	.A1(dataIn[9]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U304 (
	.ZN(\regIn[27][8] ),
	.A(n224), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U305 (
	.ZN(n224),
	.B2(\regOut[27][8] ),
	.B1(n223),
	.A2(N366),
	.A1(dataIn[8]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U306 (
	.ZN(\regIn[27][7] ),
	.A(n225), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U307 (
	.ZN(n225),
	.B2(\regOut[27][7] ),
	.B1(n223),
	.A2(N366),
	.A1(dataIn[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U308 (
	.ZN(\regIn[27][6] ),
	.A(n226), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U309 (
	.ZN(n226),
	.B2(\regOut[27][6] ),
	.B1(n223),
	.A2(N366),
	.A1(dataIn[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U310 (
	.ZN(\regIn[27][5] ),
	.A(n227), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U311 (
	.ZN(n227),
	.B2(\regOut[27][5] ),
	.B1(n223),
	.A2(N366),
	.A1(dataIn[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U312 (
	.ZN(\regIn[27][4] ),
	.A(n228), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U313 (
	.ZN(n228),
	.B2(\regOut[27][4] ),
	.B1(n223),
	.A2(N366),
	.A1(dataIn[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U314 (
	.ZN(\regIn[27][3] ),
	.A(n229), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U315 (
	.ZN(n229),
	.B2(\regOut[27][3] ),
	.B1(n223),
	.A2(N366),
	.A1(dataIn[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U316 (
	.ZN(\regIn[27][2] ),
	.A(n230), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U317 (
	.ZN(n230),
	.B2(\regOut[27][2] ),
	.B1(n223),
	.A2(N366),
	.A1(dataIn[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U318 (
	.ZN(\regIn[27][1] ),
	.A(n231), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U319 (
	.ZN(n231),
	.B2(\regOut[27][1] ),
	.B1(n223),
	.A2(N366),
	.A1(dataIn[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U320 (
	.ZN(\regIn[27][15] ),
	.A(n232), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U321 (
	.ZN(n232),
	.B2(\regOut[27][15] ),
	.B1(n223),
	.A2(N366),
	.A1(dataIn[15]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U322 (
	.ZN(\regIn[27][14] ),
	.A(n233), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U323 (
	.ZN(n233),
	.B2(\regOut[27][14] ),
	.B1(n223),
	.A2(N366),
	.A1(dataIn[14]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U324 (
	.ZN(\regIn[27][13] ),
	.A(n234), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U325 (
	.ZN(n234),
	.B2(\regOut[27][13] ),
	.B1(n223),
	.A2(N366),
	.A1(dataIn[13]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U326 (
	.ZN(\regIn[27][12] ),
	.A(n235), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U327 (
	.ZN(n235),
	.B2(\regOut[27][12] ),
	.B1(n223),
	.A2(N366),
	.A1(dataIn[12]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U328 (
	.ZN(\regIn[27][11] ),
	.A(n236), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U329 (
	.ZN(n236),
	.B2(\regOut[27][11] ),
	.B1(n223),
	.A2(N366),
	.A1(dataIn[11]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U330 (
	.ZN(\regIn[27][10] ),
	.A(n237), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U331 (
	.ZN(n237),
	.B2(\regOut[27][10] ),
	.B1(n223),
	.A2(N366),
	.A1(dataIn[10]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U332 (
	.ZN(\regIn[27][0] ),
	.A(n238), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U333 (
	.ZN(n238),
	.B2(\regOut[27][0] ),
	.B1(n223),
	.A2(N366),
	.A1(dataIn[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U334 (
	.ZN(n223),
	.A(N366), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U335 (
	.ZN(\regIn[26][9] ),
	.A(n239), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U336 (
	.ZN(n239),
	.B2(\regOut[26][9] ),
	.B1(n240),
	.A2(N360),
	.A1(dataIn[9]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U337 (
	.ZN(\regIn[26][8] ),
	.A(n241), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U338 (
	.ZN(n241),
	.B2(\regOut[26][8] ),
	.B1(n240),
	.A2(N360),
	.A1(dataIn[8]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U339 (
	.ZN(\regIn[26][7] ),
	.A(n242), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U340 (
	.ZN(n242),
	.B2(\regOut[26][7] ),
	.B1(n240),
	.A2(N360),
	.A1(dataIn[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U341 (
	.ZN(\regIn[26][6] ),
	.A(n243), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U342 (
	.ZN(n243),
	.B2(\regOut[26][6] ),
	.B1(n240),
	.A2(N360),
	.A1(dataIn[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U343 (
	.ZN(\regIn[26][5] ),
	.A(n244), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U344 (
	.ZN(n244),
	.B2(\regOut[26][5] ),
	.B1(n240),
	.A2(N360),
	.A1(dataIn[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U345 (
	.ZN(\regIn[26][4] ),
	.A(n245), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U346 (
	.ZN(n245),
	.B2(\regOut[26][4] ),
	.B1(n240),
	.A2(N360),
	.A1(dataIn[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U347 (
	.ZN(\regIn[26][3] ),
	.A(n246), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U348 (
	.ZN(n246),
	.B2(\regOut[26][3] ),
	.B1(n240),
	.A2(N360),
	.A1(dataIn[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U349 (
	.ZN(\regIn[26][2] ),
	.A(n247), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U350 (
	.ZN(n247),
	.B2(\regOut[26][2] ),
	.B1(n240),
	.A2(N360),
	.A1(dataIn[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U351 (
	.ZN(\regIn[26][1] ),
	.A(n248), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U352 (
	.ZN(n248),
	.B2(\regOut[26][1] ),
	.B1(n240),
	.A2(N360),
	.A1(dataIn[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U353 (
	.ZN(\regIn[26][15] ),
	.A(n249), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U354 (
	.ZN(n249),
	.B2(\regOut[26][15] ),
	.B1(n240),
	.A2(N360),
	.A1(dataIn[15]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U355 (
	.ZN(\regIn[26][14] ),
	.A(n250), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U356 (
	.ZN(n250),
	.B2(\regOut[26][14] ),
	.B1(n240),
	.A2(N360),
	.A1(dataIn[14]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U357 (
	.ZN(\regIn[26][13] ),
	.A(n251), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U358 (
	.ZN(n251),
	.B2(\regOut[26][13] ),
	.B1(n240),
	.A2(N360),
	.A1(dataIn[13]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U359 (
	.ZN(\regIn[26][12] ),
	.A(n252), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U360 (
	.ZN(n252),
	.B2(\regOut[26][12] ),
	.B1(n240),
	.A2(N360),
	.A1(dataIn[12]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U361 (
	.ZN(\regIn[26][11] ),
	.A(n253), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U362 (
	.ZN(n253),
	.B2(\regOut[26][11] ),
	.B1(n240),
	.A2(N360),
	.A1(dataIn[11]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U363 (
	.ZN(\regIn[26][10] ),
	.A(n254), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U364 (
	.ZN(n254),
	.B2(\regOut[26][10] ),
	.B1(n240),
	.A2(N360),
	.A1(dataIn[10]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U365 (
	.ZN(\regIn[26][0] ),
	.A(n255), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U366 (
	.ZN(n255),
	.B2(\regOut[26][0] ),
	.B1(n240),
	.A2(N360),
	.A1(dataIn[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U367 (
	.ZN(n240),
	.A(N360), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U368 (
	.ZN(\regIn[25][9] ),
	.B2(n257),
	.B1(N354),
	.A2(n256),
	.A1(n3), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U369 (
	.ZN(\regIn[25][8] ),
	.B2(n258),
	.B1(N354),
	.A2(n256),
	.A1(n5), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U370 (
	.ZN(\regIn[25][7] ),
	.B2(n259),
	.B1(N354),
	.A2(n256),
	.A1(n7), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U371 (
	.ZN(\regIn[25][6] ),
	.B2(n260),
	.B1(N354),
	.A2(n256),
	.A1(n9), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U372 (
	.ZN(\regIn[25][5] ),
	.B2(n261),
	.B1(N354),
	.A2(n256),
	.A1(n11), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U373 (
	.ZN(\regIn[25][4] ),
	.B2(n262),
	.B1(N354),
	.A2(n256),
	.A1(n13), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U374 (
	.ZN(\regIn[25][3] ),
	.B2(n263),
	.B1(N354),
	.A2(n256),
	.A1(n15), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U375 (
	.ZN(\regIn[25][2] ),
	.B2(n264),
	.B1(N354),
	.A2(n256),
	.A1(n17), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U376 (
	.ZN(\regIn[25][1] ),
	.B2(n265),
	.B1(N354),
	.A2(n256),
	.A1(n19), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U377 (
	.ZN(\regIn[25][15] ),
	.B2(n266),
	.B1(N354),
	.A2(n256),
	.A1(n21), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U378 (
	.ZN(\regIn[25][14] ),
	.B2(n267),
	.B1(N354),
	.A2(n256),
	.A1(n23), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U379 (
	.ZN(\regIn[25][13] ),
	.B2(n268),
	.B1(N354),
	.A2(n256),
	.A1(n25), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U380 (
	.ZN(\regIn[25][12] ),
	.B2(n269),
	.B1(N354),
	.A2(n256),
	.A1(n27), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U381 (
	.ZN(\regIn[25][11] ),
	.B2(n270),
	.B1(N354),
	.A2(n256),
	.A1(n29), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U382 (
	.ZN(\regIn[25][10] ),
	.B2(n271),
	.B1(N354),
	.A2(n256),
	.A1(n31), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U383 (
	.ZN(\regIn[25][0] ),
	.B2(n272),
	.B1(N354),
	.A2(n256),
	.A1(n33), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U384 (
	.ZN(n256),
	.A(N354), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U385 (
	.ZN(\regIn[24][9] ),
	.B2(n274),
	.B1(N348),
	.A2(n273),
	.A1(n3), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U386 (
	.ZN(\regIn[24][8] ),
	.B2(n275),
	.B1(N348),
	.A2(n273),
	.A1(n5), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U387 (
	.ZN(\regIn[24][7] ),
	.B2(n276),
	.B1(N348),
	.A2(n273),
	.A1(n7), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U388 (
	.ZN(\regIn[24][6] ),
	.B2(n277),
	.B1(N348),
	.A2(n273),
	.A1(n9), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U389 (
	.ZN(\regIn[24][5] ),
	.B2(n278),
	.B1(N348),
	.A2(n273),
	.A1(n11), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U390 (
	.ZN(\regIn[24][4] ),
	.B2(n279),
	.B1(N348),
	.A2(n273),
	.A1(n13), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U391 (
	.ZN(\regIn[24][3] ),
	.B2(n280),
	.B1(N348),
	.A2(n273),
	.A1(n15), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U392 (
	.ZN(\regIn[24][2] ),
	.B2(n281),
	.B1(N348),
	.A2(n273),
	.A1(n17), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U393 (
	.ZN(\regIn[24][1] ),
	.B2(n282),
	.B1(N348),
	.A2(n273),
	.A1(n19), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U394 (
	.ZN(\regIn[24][15] ),
	.B2(n283),
	.B1(N348),
	.A2(n273),
	.A1(n21), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U395 (
	.ZN(\regIn[24][14] ),
	.B2(n284),
	.B1(N348),
	.A2(n273),
	.A1(n23), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U396 (
	.ZN(\regIn[24][13] ),
	.B2(n285),
	.B1(N348),
	.A2(n273),
	.A1(n25), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U397 (
	.ZN(\regIn[24][12] ),
	.B2(n286),
	.B1(N348),
	.A2(n273),
	.A1(n27), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U398 (
	.ZN(\regIn[24][11] ),
	.B2(n287),
	.B1(N348),
	.A2(n273),
	.A1(n29), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U399 (
	.ZN(\regIn[24][10] ),
	.B2(n288),
	.B1(N348),
	.A2(n273),
	.A1(n31), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U400 (
	.ZN(\regIn[24][0] ),
	.B2(n289),
	.B1(N348),
	.A2(n273),
	.A1(n33), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U401 (
	.ZN(n273),
	.A(N348), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U402 (
	.ZN(\regIn[23][9] ),
	.A(n290), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U403 (
	.ZN(n290),
	.B2(\regOut[23][9] ),
	.B1(n291),
	.A2(N342),
	.A1(dataIn[9]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U404 (
	.ZN(\regIn[23][8] ),
	.A(n292), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U405 (
	.ZN(n292),
	.B2(\regOut[23][8] ),
	.B1(n291),
	.A2(N342),
	.A1(dataIn[8]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U406 (
	.ZN(\regIn[23][7] ),
	.A(n293), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U407 (
	.ZN(n293),
	.B2(\regOut[23][7] ),
	.B1(n291),
	.A2(N342),
	.A1(dataIn[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U408 (
	.ZN(\regIn[23][6] ),
	.A(n294), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U409 (
	.ZN(n294),
	.B2(\regOut[23][6] ),
	.B1(n291),
	.A2(N342),
	.A1(dataIn[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U410 (
	.ZN(\regIn[23][5] ),
	.A(n295), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U411 (
	.ZN(n295),
	.B2(\regOut[23][5] ),
	.B1(n291),
	.A2(N342),
	.A1(dataIn[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U412 (
	.ZN(\regIn[23][4] ),
	.A(n296), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U413 (
	.ZN(n296),
	.B2(\regOut[23][4] ),
	.B1(n291),
	.A2(N342),
	.A1(dataIn[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U414 (
	.ZN(\regIn[23][3] ),
	.A(n297), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U415 (
	.ZN(n297),
	.B2(\regOut[23][3] ),
	.B1(n291),
	.A2(N342),
	.A1(dataIn[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U416 (
	.ZN(\regIn[23][2] ),
	.A(n298), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U417 (
	.ZN(n298),
	.B2(\regOut[23][2] ),
	.B1(n291),
	.A2(N342),
	.A1(dataIn[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U418 (
	.ZN(\regIn[23][1] ),
	.A(n299), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U419 (
	.ZN(n299),
	.B2(\regOut[23][1] ),
	.B1(n291),
	.A2(N342),
	.A1(dataIn[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U420 (
	.ZN(\regIn[23][15] ),
	.A(n300), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U421 (
	.ZN(n300),
	.B2(\regOut[23][15] ),
	.B1(n291),
	.A2(N342),
	.A1(dataIn[15]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U422 (
	.ZN(\regIn[23][14] ),
	.A(n301), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U423 (
	.ZN(n301),
	.B2(\regOut[23][14] ),
	.B1(n291),
	.A2(N342),
	.A1(dataIn[14]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U424 (
	.ZN(\regIn[23][13] ),
	.A(n302), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U425 (
	.ZN(n302),
	.B2(\regOut[23][13] ),
	.B1(n291),
	.A2(N342),
	.A1(dataIn[13]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U426 (
	.ZN(\regIn[23][12] ),
	.A(n303), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U427 (
	.ZN(n303),
	.B2(\regOut[23][12] ),
	.B1(n291),
	.A2(N342),
	.A1(dataIn[12]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U428 (
	.ZN(\regIn[23][11] ),
	.A(n304), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U429 (
	.ZN(n304),
	.B2(\regOut[23][11] ),
	.B1(n291),
	.A2(N342),
	.A1(dataIn[11]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U430 (
	.ZN(\regIn[23][10] ),
	.A(n305), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U431 (
	.ZN(n305),
	.B2(\regOut[23][10] ),
	.B1(n291),
	.A2(N342),
	.A1(dataIn[10]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U432 (
	.ZN(\regIn[23][0] ),
	.A(n306), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U433 (
	.ZN(n306),
	.B2(\regOut[23][0] ),
	.B1(n291),
	.A2(N342),
	.A1(dataIn[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U434 (
	.ZN(n291),
	.A(N342), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U435 (
	.ZN(\regIn[22][9] ),
	.A(n307), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U436 (
	.ZN(n307),
	.B2(\regOut[22][9] ),
	.B1(n308),
	.A2(N336),
	.A1(dataIn[9]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U437 (
	.ZN(\regIn[22][8] ),
	.A(n309), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U438 (
	.ZN(n309),
	.B2(\regOut[22][8] ),
	.B1(n308),
	.A2(N336),
	.A1(dataIn[8]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U439 (
	.ZN(\regIn[22][7] ),
	.A(n310), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U440 (
	.ZN(n310),
	.B2(\regOut[22][7] ),
	.B1(n308),
	.A2(N336),
	.A1(dataIn[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U441 (
	.ZN(\regIn[22][6] ),
	.A(n311), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U442 (
	.ZN(n311),
	.B2(\regOut[22][6] ),
	.B1(n308),
	.A2(N336),
	.A1(dataIn[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U443 (
	.ZN(\regIn[22][5] ),
	.A(n312), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U444 (
	.ZN(n312),
	.B2(\regOut[22][5] ),
	.B1(n308),
	.A2(N336),
	.A1(dataIn[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U445 (
	.ZN(\regIn[22][4] ),
	.A(n313), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U446 (
	.ZN(n313),
	.B2(\regOut[22][4] ),
	.B1(n308),
	.A2(N336),
	.A1(dataIn[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U447 (
	.ZN(\regIn[22][3] ),
	.A(n314), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U448 (
	.ZN(n314),
	.B2(\regOut[22][3] ),
	.B1(n308),
	.A2(N336),
	.A1(dataIn[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U449 (
	.ZN(\regIn[22][2] ),
	.A(n315), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U450 (
	.ZN(n315),
	.B2(\regOut[22][2] ),
	.B1(n308),
	.A2(N336),
	.A1(dataIn[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U451 (
	.ZN(\regIn[22][1] ),
	.A(n316), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U452 (
	.ZN(n316),
	.B2(\regOut[22][1] ),
	.B1(n308),
	.A2(N336),
	.A1(dataIn[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U453 (
	.ZN(\regIn[22][15] ),
	.A(n317), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U454 (
	.ZN(n317),
	.B2(\regOut[22][15] ),
	.B1(n308),
	.A2(N336),
	.A1(dataIn[15]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U455 (
	.ZN(\regIn[22][14] ),
	.A(n318), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U456 (
	.ZN(n318),
	.B2(\regOut[22][14] ),
	.B1(n308),
	.A2(N336),
	.A1(dataIn[14]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U457 (
	.ZN(\regIn[22][13] ),
	.A(n319), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U458 (
	.ZN(n319),
	.B2(\regOut[22][13] ),
	.B1(n308),
	.A2(N336),
	.A1(dataIn[13]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U459 (
	.ZN(\regIn[22][12] ),
	.A(n320), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U460 (
	.ZN(n320),
	.B2(\regOut[22][12] ),
	.B1(n308),
	.A2(N336),
	.A1(dataIn[12]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U461 (
	.ZN(\regIn[22][11] ),
	.A(n321), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U462 (
	.ZN(n321),
	.B2(\regOut[22][11] ),
	.B1(n308),
	.A2(N336),
	.A1(dataIn[11]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U463 (
	.ZN(\regIn[22][10] ),
	.A(n322), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U464 (
	.ZN(n322),
	.B2(\regOut[22][10] ),
	.B1(n308),
	.A2(N336),
	.A1(dataIn[10]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U465 (
	.ZN(\regIn[22][0] ),
	.A(n323), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U466 (
	.ZN(n323),
	.B2(\regOut[22][0] ),
	.B1(n308),
	.A2(N336),
	.A1(dataIn[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U467 (
	.ZN(n308),
	.A(N336), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U468 (
	.ZN(\regIn[21][9] ),
	.B2(n325),
	.B1(N330),
	.A2(n324),
	.A1(n3), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U469 (
	.ZN(\regIn[21][8] ),
	.B2(n326),
	.B1(N330),
	.A2(n324),
	.A1(n5), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U470 (
	.ZN(\regIn[21][7] ),
	.B2(n327),
	.B1(N330),
	.A2(n324),
	.A1(n7), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U471 (
	.ZN(\regIn[21][6] ),
	.B2(n328),
	.B1(N330),
	.A2(n324),
	.A1(n9), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U472 (
	.ZN(\regIn[21][5] ),
	.B2(n329),
	.B1(N330),
	.A2(n324),
	.A1(n11), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U473 (
	.ZN(\regIn[21][4] ),
	.B2(n330),
	.B1(N330),
	.A2(n324),
	.A1(n13), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U474 (
	.ZN(\regIn[21][3] ),
	.B2(n331),
	.B1(N330),
	.A2(n324),
	.A1(n15), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U475 (
	.ZN(\regIn[21][2] ),
	.B2(n332),
	.B1(N330),
	.A2(n324),
	.A1(n17), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U476 (
	.ZN(\regIn[21][1] ),
	.B2(n333),
	.B1(N330),
	.A2(n324),
	.A1(n19), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U477 (
	.ZN(\regIn[21][15] ),
	.B2(n334),
	.B1(N330),
	.A2(n324),
	.A1(n21), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U478 (
	.ZN(\regIn[21][14] ),
	.B2(n335),
	.B1(N330),
	.A2(n324),
	.A1(n23), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U479 (
	.ZN(\regIn[21][13] ),
	.B2(n336),
	.B1(N330),
	.A2(n324),
	.A1(n25), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U480 (
	.ZN(\regIn[21][12] ),
	.B2(n337),
	.B1(N330),
	.A2(n324),
	.A1(n27), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U481 (
	.ZN(\regIn[21][11] ),
	.B2(n338),
	.B1(N330),
	.A2(n324),
	.A1(n29), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U482 (
	.ZN(\regIn[21][10] ),
	.B2(n339),
	.B1(N330),
	.A2(n324),
	.A1(n31), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U483 (
	.ZN(\regIn[21][0] ),
	.B2(n340),
	.B1(N330),
	.A2(n324),
	.A1(n33), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U484 (
	.ZN(n324),
	.A(N330), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U485 (
	.ZN(\regIn[20][9] ),
	.B2(n342),
	.B1(N324),
	.A2(n341),
	.A1(n3), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U486 (
	.ZN(\regIn[20][8] ),
	.B2(n343),
	.B1(N324),
	.A2(n341),
	.A1(n5), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U487 (
	.ZN(\regIn[20][7] ),
	.B2(n344),
	.B1(N324),
	.A2(n341),
	.A1(n7), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U488 (
	.ZN(\regIn[20][6] ),
	.B2(n345),
	.B1(N324),
	.A2(n341),
	.A1(n9), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U489 (
	.ZN(\regIn[20][5] ),
	.B2(n346),
	.B1(N324),
	.A2(n341),
	.A1(n11), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U490 (
	.ZN(\regIn[20][4] ),
	.B2(n347),
	.B1(N324),
	.A2(n341),
	.A1(n13), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U491 (
	.ZN(\regIn[20][3] ),
	.B2(n348),
	.B1(N324),
	.A2(n341),
	.A1(n15), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U492 (
	.ZN(\regIn[20][2] ),
	.B2(n349),
	.B1(N324),
	.A2(n341),
	.A1(n17), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U493 (
	.ZN(\regIn[20][1] ),
	.B2(n350),
	.B1(N324),
	.A2(n341),
	.A1(n19), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U494 (
	.ZN(\regIn[20][15] ),
	.B2(n351),
	.B1(N324),
	.A2(n341),
	.A1(n21), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U495 (
	.ZN(\regIn[20][14] ),
	.B2(n352),
	.B1(N324),
	.A2(n341),
	.A1(n23), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U496 (
	.ZN(\regIn[20][13] ),
	.B2(n353),
	.B1(N324),
	.A2(n341),
	.A1(n25), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U497 (
	.ZN(\regIn[20][12] ),
	.B2(n354),
	.B1(N324),
	.A2(n341),
	.A1(n27), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U498 (
	.ZN(\regIn[20][11] ),
	.B2(n355),
	.B1(N324),
	.A2(n341),
	.A1(n29), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U499 (
	.ZN(\regIn[20][10] ),
	.B2(n356),
	.B1(N324),
	.A2(n341),
	.A1(n31), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U500 (
	.ZN(\regIn[20][0] ),
	.B2(n357),
	.B1(N324),
	.A2(n341),
	.A1(n33), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U501 (
	.ZN(n341),
	.A(N324), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U502 (
	.ZN(\regIn[1][9] ),
	.B2(n359),
	.B1(N206),
	.A2(n358),
	.A1(n3), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U503 (
	.ZN(\regIn[1][8] ),
	.B2(n360),
	.B1(N206),
	.A2(n358),
	.A1(n5), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U504 (
	.ZN(\regIn[1][7] ),
	.B2(n361),
	.B1(N206),
	.A2(n358),
	.A1(n7), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U505 (
	.ZN(\regIn[1][6] ),
	.B2(n362),
	.B1(N206),
	.A2(n358),
	.A1(n9), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U506 (
	.ZN(\regIn[1][5] ),
	.B2(n363),
	.B1(N206),
	.A2(n358),
	.A1(n11), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U507 (
	.ZN(\regIn[1][4] ),
	.B2(n364),
	.B1(N206),
	.A2(n358),
	.A1(n13), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U508 (
	.ZN(\regIn[1][3] ),
	.B2(n365),
	.B1(N206),
	.A2(n358),
	.A1(n15), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U509 (
	.ZN(\regIn[1][2] ),
	.B2(n366),
	.B1(N206),
	.A2(n358),
	.A1(n17), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U510 (
	.ZN(\regIn[1][1] ),
	.B2(n367),
	.B1(N206),
	.A2(n358),
	.A1(n19), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U511 (
	.ZN(\regIn[1][15] ),
	.B2(n368),
	.B1(N206),
	.A2(n358),
	.A1(n21), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U512 (
	.ZN(\regIn[1][14] ),
	.B2(n369),
	.B1(N206),
	.A2(n358),
	.A1(n23), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U513 (
	.ZN(\regIn[1][13] ),
	.B2(n370),
	.B1(N206),
	.A2(n358),
	.A1(n25), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U514 (
	.ZN(\regIn[1][12] ),
	.B2(n371),
	.B1(N206),
	.A2(n358),
	.A1(n27), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U515 (
	.ZN(\regIn[1][11] ),
	.B2(n372),
	.B1(N206),
	.A2(n358),
	.A1(n29), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U516 (
	.ZN(\regIn[1][10] ),
	.B2(n373),
	.B1(N206),
	.A2(n358),
	.A1(n31), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U517 (
	.ZN(\regIn[1][0] ),
	.B2(n374),
	.B1(N206),
	.A2(n358),
	.A1(n33), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U518 (
	.ZN(n358),
	.A(N206), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U519 (
	.ZN(\regIn[19][9] ),
	.A(n375), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U520 (
	.ZN(n375),
	.B2(\regOut[19][9] ),
	.B1(n376),
	.A2(N318),
	.A1(dataIn[9]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U521 (
	.ZN(\regIn[19][8] ),
	.A(n377), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U522 (
	.ZN(n377),
	.B2(\regOut[19][8] ),
	.B1(n376),
	.A2(N318),
	.A1(dataIn[8]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U523 (
	.ZN(\regIn[19][7] ),
	.A(n378), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U524 (
	.ZN(n378),
	.B2(\regOut[19][7] ),
	.B1(n376),
	.A2(N318),
	.A1(dataIn[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U525 (
	.ZN(\regIn[19][6] ),
	.A(n379), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U526 (
	.ZN(n379),
	.B2(\regOut[19][6] ),
	.B1(n376),
	.A2(N318),
	.A1(dataIn[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U527 (
	.ZN(\regIn[19][5] ),
	.A(n380), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U528 (
	.ZN(n380),
	.B2(\regOut[19][5] ),
	.B1(n376),
	.A2(N318),
	.A1(dataIn[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U529 (
	.ZN(\regIn[19][4] ),
	.A(n381), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U530 (
	.ZN(n381),
	.B2(\regOut[19][4] ),
	.B1(n376),
	.A2(N318),
	.A1(dataIn[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U531 (
	.ZN(\regIn[19][3] ),
	.A(n382), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U532 (
	.ZN(n382),
	.B2(\regOut[19][3] ),
	.B1(n376),
	.A2(N318),
	.A1(dataIn[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U533 (
	.ZN(\regIn[19][2] ),
	.A(n383), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U534 (
	.ZN(n383),
	.B2(\regOut[19][2] ),
	.B1(n376),
	.A2(N318),
	.A1(dataIn[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U535 (
	.ZN(\regIn[19][1] ),
	.A(n384), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U536 (
	.ZN(n384),
	.B2(\regOut[19][1] ),
	.B1(n376),
	.A2(N318),
	.A1(dataIn[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U537 (
	.ZN(\regIn[19][15] ),
	.A(n385), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U538 (
	.ZN(n385),
	.B2(\regOut[19][15] ),
	.B1(n376),
	.A2(N318),
	.A1(dataIn[15]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U539 (
	.ZN(\regIn[19][14] ),
	.A(n386), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U540 (
	.ZN(n386),
	.B2(\regOut[19][14] ),
	.B1(n376),
	.A2(N318),
	.A1(dataIn[14]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U541 (
	.ZN(\regIn[19][13] ),
	.A(n387), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U542 (
	.ZN(n387),
	.B2(\regOut[19][13] ),
	.B1(n376),
	.A2(N318),
	.A1(dataIn[13]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U543 (
	.ZN(\regIn[19][12] ),
	.A(n388), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U544 (
	.ZN(n388),
	.B2(\regOut[19][12] ),
	.B1(n376),
	.A2(N318),
	.A1(dataIn[12]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U545 (
	.ZN(\regIn[19][11] ),
	.A(n389), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U546 (
	.ZN(n389),
	.B2(\regOut[19][11] ),
	.B1(n376),
	.A2(N318),
	.A1(dataIn[11]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U547 (
	.ZN(\regIn[19][10] ),
	.A(n390), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U548 (
	.ZN(n390),
	.B2(\regOut[19][10] ),
	.B1(n376),
	.A2(N318),
	.A1(dataIn[10]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U549 (
	.ZN(\regIn[19][0] ),
	.A(n391), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U550 (
	.ZN(n391),
	.B2(\regOut[19][0] ),
	.B1(n376),
	.A2(N318),
	.A1(dataIn[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U551 (
	.ZN(n376),
	.A(N318), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U552 (
	.ZN(\regIn[18][9] ),
	.A(n392), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U553 (
	.ZN(n392),
	.B2(\regOut[18][9] ),
	.B1(n393),
	.A2(N312),
	.A1(dataIn[9]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U554 (
	.ZN(\regIn[18][8] ),
	.A(n394), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U555 (
	.ZN(n394),
	.B2(\regOut[18][8] ),
	.B1(n393),
	.A2(N312),
	.A1(dataIn[8]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U556 (
	.ZN(\regIn[18][7] ),
	.A(n395), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U557 (
	.ZN(n395),
	.B2(\regOut[18][7] ),
	.B1(n393),
	.A2(N312),
	.A1(dataIn[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U558 (
	.ZN(\regIn[18][6] ),
	.A(n396), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U559 (
	.ZN(n396),
	.B2(\regOut[18][6] ),
	.B1(n393),
	.A2(N312),
	.A1(dataIn[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U560 (
	.ZN(\regIn[18][5] ),
	.A(n397), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U561 (
	.ZN(n397),
	.B2(\regOut[18][5] ),
	.B1(n393),
	.A2(N312),
	.A1(dataIn[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U562 (
	.ZN(\regIn[18][4] ),
	.A(n398), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U563 (
	.ZN(n398),
	.B2(\regOut[18][4] ),
	.B1(n393),
	.A2(N312),
	.A1(dataIn[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U564 (
	.ZN(\regIn[18][3] ),
	.A(n399), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U565 (
	.ZN(n399),
	.B2(\regOut[18][3] ),
	.B1(n393),
	.A2(N312),
	.A1(dataIn[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U566 (
	.ZN(\regIn[18][2] ),
	.A(n400), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U567 (
	.ZN(n400),
	.B2(\regOut[18][2] ),
	.B1(n393),
	.A2(N312),
	.A1(dataIn[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U568 (
	.ZN(\regIn[18][1] ),
	.A(n401), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U569 (
	.ZN(n401),
	.B2(\regOut[18][1] ),
	.B1(n393),
	.A2(N312),
	.A1(dataIn[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U570 (
	.ZN(\regIn[18][15] ),
	.A(n402), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U571 (
	.ZN(n402),
	.B2(\regOut[18][15] ),
	.B1(n393),
	.A2(N312),
	.A1(dataIn[15]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U572 (
	.ZN(\regIn[18][14] ),
	.A(n403), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U573 (
	.ZN(n403),
	.B2(\regOut[18][14] ),
	.B1(n393),
	.A2(N312),
	.A1(dataIn[14]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U574 (
	.ZN(\regIn[18][13] ),
	.A(n404), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U575 (
	.ZN(n404),
	.B2(\regOut[18][13] ),
	.B1(n393),
	.A2(N312),
	.A1(dataIn[13]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U576 (
	.ZN(\regIn[18][12] ),
	.A(n405), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U577 (
	.ZN(n405),
	.B2(\regOut[18][12] ),
	.B1(n393),
	.A2(N312),
	.A1(dataIn[12]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U578 (
	.ZN(\regIn[18][11] ),
	.A(n406), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U579 (
	.ZN(n406),
	.B2(\regOut[18][11] ),
	.B1(n393),
	.A2(N312),
	.A1(dataIn[11]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U580 (
	.ZN(\regIn[18][10] ),
	.A(n407), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U581 (
	.ZN(n407),
	.B2(\regOut[18][10] ),
	.B1(n393),
	.A2(N312),
	.A1(dataIn[10]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U582 (
	.ZN(\regIn[18][0] ),
	.A(n408), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U583 (
	.ZN(n408),
	.B2(\regOut[18][0] ),
	.B1(n393),
	.A2(N312),
	.A1(dataIn[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U584 (
	.ZN(n393),
	.A(N312), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U585 (
	.ZN(\regIn[17][9] ),
	.B2(n410),
	.B1(N306),
	.A2(n409),
	.A1(n3), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U586 (
	.ZN(\regIn[17][8] ),
	.B2(n411),
	.B1(N306),
	.A2(n409),
	.A1(n5), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U587 (
	.ZN(\regIn[17][7] ),
	.B2(n412),
	.B1(N306),
	.A2(n409),
	.A1(n7), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U588 (
	.ZN(\regIn[17][6] ),
	.B2(n413),
	.B1(N306),
	.A2(n409),
	.A1(n9), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U589 (
	.ZN(\regIn[17][5] ),
	.B2(n414),
	.B1(N306),
	.A2(n409),
	.A1(n11), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U590 (
	.ZN(\regIn[17][4] ),
	.B2(n415),
	.B1(N306),
	.A2(n409),
	.A1(n13), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U591 (
	.ZN(\regIn[17][3] ),
	.B2(n416),
	.B1(N306),
	.A2(n409),
	.A1(n15), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U592 (
	.ZN(\regIn[17][2] ),
	.B2(n417),
	.B1(N306),
	.A2(n409),
	.A1(n17), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U593 (
	.ZN(\regIn[17][1] ),
	.B2(n418),
	.B1(N306),
	.A2(n409),
	.A1(n19), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U594 (
	.ZN(\regIn[17][15] ),
	.B2(n419),
	.B1(N306),
	.A2(n409),
	.A1(n21), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U595 (
	.ZN(\regIn[17][14] ),
	.B2(n420),
	.B1(N306),
	.A2(n409),
	.A1(n23), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U596 (
	.ZN(\regIn[17][13] ),
	.B2(n421),
	.B1(N306),
	.A2(n409),
	.A1(n25), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U597 (
	.ZN(\regIn[17][12] ),
	.B2(n422),
	.B1(N306),
	.A2(n409),
	.A1(n27), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U598 (
	.ZN(\regIn[17][11] ),
	.B2(n423),
	.B1(N306),
	.A2(n409),
	.A1(n29), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U599 (
	.ZN(\regIn[17][10] ),
	.B2(n424),
	.B1(N306),
	.A2(n409),
	.A1(n31), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U600 (
	.ZN(\regIn[17][0] ),
	.B2(n425),
	.B1(N306),
	.A2(n409),
	.A1(n33), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U601 (
	.ZN(n409),
	.A(N306), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U602 (
	.ZN(\regIn[16][9] ),
	.B2(n427),
	.B1(N300),
	.A2(n426),
	.A1(n3), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U603 (
	.ZN(\regIn[16][8] ),
	.B2(n428),
	.B1(N300),
	.A2(n426),
	.A1(n5), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U604 (
	.ZN(\regIn[16][7] ),
	.B2(n429),
	.B1(N300),
	.A2(n426),
	.A1(n7), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U605 (
	.ZN(\regIn[16][6] ),
	.B2(n430),
	.B1(N300),
	.A2(n426),
	.A1(n9), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U606 (
	.ZN(\regIn[16][5] ),
	.B2(n431),
	.B1(N300),
	.A2(n426),
	.A1(n11), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U607 (
	.ZN(\regIn[16][4] ),
	.B2(n432),
	.B1(N300),
	.A2(n426),
	.A1(n13), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U608 (
	.ZN(\regIn[16][3] ),
	.B2(n433),
	.B1(N300),
	.A2(n426),
	.A1(n15), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U609 (
	.ZN(\regIn[16][2] ),
	.B2(n434),
	.B1(N300),
	.A2(n426),
	.A1(n17), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U610 (
	.ZN(\regIn[16][1] ),
	.B2(n435),
	.B1(N300),
	.A2(n426),
	.A1(n19), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U611 (
	.ZN(\regIn[16][15] ),
	.B2(n436),
	.B1(N300),
	.A2(n426),
	.A1(n21), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U612 (
	.ZN(\regIn[16][14] ),
	.B2(n437),
	.B1(N300),
	.A2(n426),
	.A1(n23), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U613 (
	.ZN(\regIn[16][13] ),
	.B2(n438),
	.B1(N300),
	.A2(n426),
	.A1(n25), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U614 (
	.ZN(\regIn[16][12] ),
	.B2(n439),
	.B1(N300),
	.A2(n426),
	.A1(n27), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U615 (
	.ZN(\regIn[16][11] ),
	.B2(n440),
	.B1(N300),
	.A2(n426),
	.A1(n29), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U616 (
	.ZN(\regIn[16][10] ),
	.B2(n441),
	.B1(N300),
	.A2(n426),
	.A1(n31), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U617 (
	.ZN(\regIn[16][0] ),
	.B2(n442),
	.B1(N300),
	.A2(n426),
	.A1(n33), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U618 (
	.ZN(n426),
	.A(N300), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U619 (
	.ZN(\regIn[15][9] ),
	.A(n443), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U620 (
	.ZN(n443),
	.B2(\regOut[15][9] ),
	.B1(n444),
	.A2(N293),
	.A1(dataIn[9]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U621 (
	.ZN(\regIn[15][8] ),
	.A(n445), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U622 (
	.ZN(n445),
	.B2(\regOut[15][8] ),
	.B1(n444),
	.A2(N293),
	.A1(dataIn[8]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U623 (
	.ZN(\regIn[15][7] ),
	.A(n446), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U624 (
	.ZN(n446),
	.B2(\regOut[15][7] ),
	.B1(n444),
	.A2(N293),
	.A1(dataIn[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U625 (
	.ZN(\regIn[15][6] ),
	.A(n447), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U626 (
	.ZN(n447),
	.B2(\regOut[15][6] ),
	.B1(n444),
	.A2(N293),
	.A1(dataIn[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U627 (
	.ZN(\regIn[15][5] ),
	.A(n448), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U628 (
	.ZN(n448),
	.B2(\regOut[15][5] ),
	.B1(n444),
	.A2(N293),
	.A1(dataIn[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U629 (
	.ZN(\regIn[15][4] ),
	.A(n449), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U630 (
	.ZN(n449),
	.B2(\regOut[15][4] ),
	.B1(n444),
	.A2(N293),
	.A1(dataIn[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U631 (
	.ZN(\regIn[15][3] ),
	.A(n450), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U632 (
	.ZN(n450),
	.B2(\regOut[15][3] ),
	.B1(n444),
	.A2(N293),
	.A1(dataIn[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U633 (
	.ZN(\regIn[15][2] ),
	.A(n451), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U634 (
	.ZN(n451),
	.B2(\regOut[15][2] ),
	.B1(n444),
	.A2(N293),
	.A1(dataIn[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U635 (
	.ZN(\regIn[15][1] ),
	.A(n452), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U636 (
	.ZN(n452),
	.B2(\regOut[15][1] ),
	.B1(n444),
	.A2(N293),
	.A1(dataIn[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U637 (
	.ZN(\regIn[15][15] ),
	.A(n453), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U638 (
	.ZN(n453),
	.B2(\regOut[15][15] ),
	.B1(n444),
	.A2(N293),
	.A1(dataIn[15]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U639 (
	.ZN(\regIn[15][14] ),
	.A(n454), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U640 (
	.ZN(n454),
	.B2(\regOut[15][14] ),
	.B1(n444),
	.A2(N293),
	.A1(dataIn[14]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U641 (
	.ZN(\regIn[15][13] ),
	.A(n455), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U642 (
	.ZN(n455),
	.B2(\regOut[15][13] ),
	.B1(n444),
	.A2(N293),
	.A1(dataIn[13]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U643 (
	.ZN(\regIn[15][12] ),
	.A(n456), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U644 (
	.ZN(n456),
	.B2(\regOut[15][12] ),
	.B1(n444),
	.A2(N293),
	.A1(dataIn[12]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U645 (
	.ZN(\regIn[15][11] ),
	.A(n457), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U646 (
	.ZN(n457),
	.B2(\regOut[15][11] ),
	.B1(n444),
	.A2(N293),
	.A1(dataIn[11]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U647 (
	.ZN(\regIn[15][10] ),
	.A(n458), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U648 (
	.ZN(n458),
	.B2(\regOut[15][10] ),
	.B1(n444),
	.A2(N293),
	.A1(dataIn[10]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U649 (
	.ZN(\regIn[15][0] ),
	.A(n459), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U650 (
	.ZN(n459),
	.B2(\regOut[15][0] ),
	.B1(n444),
	.A2(N293),
	.A1(dataIn[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U651 (
	.ZN(n444),
	.A(N293), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U652 (
	.ZN(\regIn[14][9] ),
	.A(n460), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U653 (
	.ZN(n460),
	.B2(\regOut[14][9] ),
	.B1(n461),
	.A2(N287),
	.A1(dataIn[9]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U654 (
	.ZN(\regIn[14][8] ),
	.A(n462), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U655 (
	.ZN(n462),
	.B2(\regOut[14][8] ),
	.B1(n461),
	.A2(N287),
	.A1(dataIn[8]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U656 (
	.ZN(\regIn[14][7] ),
	.A(n463), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U657 (
	.ZN(n463),
	.B2(\regOut[14][7] ),
	.B1(n461),
	.A2(N287),
	.A1(dataIn[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U658 (
	.ZN(\regIn[14][6] ),
	.A(n464), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U659 (
	.ZN(n464),
	.B2(\regOut[14][6] ),
	.B1(n461),
	.A2(N287),
	.A1(dataIn[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U660 (
	.ZN(\regIn[14][5] ),
	.A(n465), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U661 (
	.ZN(n465),
	.B2(\regOut[14][5] ),
	.B1(n461),
	.A2(N287),
	.A1(dataIn[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U662 (
	.ZN(\regIn[14][4] ),
	.A(n466), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U663 (
	.ZN(n466),
	.B2(\regOut[14][4] ),
	.B1(n461),
	.A2(N287),
	.A1(dataIn[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U664 (
	.ZN(\regIn[14][3] ),
	.A(n467), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U665 (
	.ZN(n467),
	.B2(\regOut[14][3] ),
	.B1(n461),
	.A2(N287),
	.A1(dataIn[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U666 (
	.ZN(\regIn[14][2] ),
	.A(n468), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U667 (
	.ZN(n468),
	.B2(\regOut[14][2] ),
	.B1(n461),
	.A2(N287),
	.A1(dataIn[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U668 (
	.ZN(\regIn[14][1] ),
	.A(n469), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U669 (
	.ZN(n469),
	.B2(\regOut[14][1] ),
	.B1(n461),
	.A2(N287),
	.A1(dataIn[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U670 (
	.ZN(\regIn[14][15] ),
	.A(n470), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U671 (
	.ZN(n470),
	.B2(\regOut[14][15] ),
	.B1(n461),
	.A2(N287),
	.A1(dataIn[15]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U672 (
	.ZN(\regIn[14][14] ),
	.A(n471), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U673 (
	.ZN(n471),
	.B2(\regOut[14][14] ),
	.B1(n461),
	.A2(N287),
	.A1(dataIn[14]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U674 (
	.ZN(\regIn[14][13] ),
	.A(n472), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U675 (
	.ZN(n472),
	.B2(\regOut[14][13] ),
	.B1(n461),
	.A2(N287),
	.A1(dataIn[13]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U676 (
	.ZN(\regIn[14][12] ),
	.A(n473), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U677 (
	.ZN(n473),
	.B2(\regOut[14][12] ),
	.B1(n461),
	.A2(N287),
	.A1(dataIn[12]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U678 (
	.ZN(\regIn[14][11] ),
	.A(n474), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U679 (
	.ZN(n474),
	.B2(\regOut[14][11] ),
	.B1(n461),
	.A2(N287),
	.A1(dataIn[11]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U680 (
	.ZN(\regIn[14][10] ),
	.A(n475), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U681 (
	.ZN(n475),
	.B2(\regOut[14][10] ),
	.B1(n461),
	.A2(N287),
	.A1(dataIn[10]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U682 (
	.ZN(\regIn[14][0] ),
	.A(n476), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U683 (
	.ZN(n476),
	.B2(\regOut[14][0] ),
	.B1(n461),
	.A2(N287),
	.A1(dataIn[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U684 (
	.ZN(n461),
	.A(N287), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U685 (
	.ZN(\regIn[13][9] ),
	.B2(n478),
	.B1(N281),
	.A2(n477),
	.A1(n3), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U686 (
	.ZN(\regIn[13][8] ),
	.B2(n479),
	.B1(N281),
	.A2(n477),
	.A1(n5), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U687 (
	.ZN(\regIn[13][7] ),
	.B2(n480),
	.B1(N281),
	.A2(n477),
	.A1(n7), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U688 (
	.ZN(\regIn[13][6] ),
	.B2(n481),
	.B1(N281),
	.A2(n477),
	.A1(n9), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U689 (
	.ZN(\regIn[13][5] ),
	.B2(n482),
	.B1(N281),
	.A2(n477),
	.A1(n11), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U690 (
	.ZN(\regIn[13][4] ),
	.B2(n483),
	.B1(N281),
	.A2(n477),
	.A1(n13), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U691 (
	.ZN(\regIn[13][3] ),
	.B2(n484),
	.B1(N281),
	.A2(n477),
	.A1(n15), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U692 (
	.ZN(\regIn[13][2] ),
	.B2(n485),
	.B1(N281),
	.A2(n477),
	.A1(n17), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U693 (
	.ZN(\regIn[13][1] ),
	.B2(n486),
	.B1(N281),
	.A2(n477),
	.A1(n19), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U694 (
	.ZN(\regIn[13][15] ),
	.B2(n487),
	.B1(N281),
	.A2(n477),
	.A1(n21), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U695 (
	.ZN(\regIn[13][14] ),
	.B2(n488),
	.B1(N281),
	.A2(n477),
	.A1(n23), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U696 (
	.ZN(\regIn[13][13] ),
	.B2(n489),
	.B1(N281),
	.A2(n477),
	.A1(n25), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U697 (
	.ZN(\regIn[13][12] ),
	.B2(n490),
	.B1(N281),
	.A2(n477),
	.A1(n27), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U698 (
	.ZN(\regIn[13][11] ),
	.B2(n491),
	.B1(N281),
	.A2(n477),
	.A1(n29), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U699 (
	.ZN(\regIn[13][10] ),
	.B2(n492),
	.B1(N281),
	.A2(n477),
	.A1(n31), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U700 (
	.ZN(\regIn[13][0] ),
	.B2(n493),
	.B1(N281),
	.A2(n477),
	.A1(n33), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U701 (
	.ZN(n477),
	.A(N281), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U702 (
	.ZN(\regIn[12][9] ),
	.B2(n495),
	.B1(N275),
	.A2(n494),
	.A1(n3), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U703 (
	.ZN(\regIn[12][8] ),
	.B2(n496),
	.B1(N275),
	.A2(n494),
	.A1(n5), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U704 (
	.ZN(\regIn[12][7] ),
	.B2(n497),
	.B1(N275),
	.A2(n494),
	.A1(n7), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U705 (
	.ZN(\regIn[12][6] ),
	.B2(n498),
	.B1(N275),
	.A2(n494),
	.A1(n9), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U706 (
	.ZN(\regIn[12][5] ),
	.B2(n499),
	.B1(N275),
	.A2(n494),
	.A1(n11), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U707 (
	.ZN(\regIn[12][4] ),
	.B2(n500),
	.B1(N275),
	.A2(n494),
	.A1(n13), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U708 (
	.ZN(\regIn[12][3] ),
	.B2(n501),
	.B1(N275),
	.A2(n494),
	.A1(n15), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U709 (
	.ZN(\regIn[12][2] ),
	.B2(n502),
	.B1(N275),
	.A2(n494),
	.A1(n17), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U710 (
	.ZN(\regIn[12][1] ),
	.B2(n503),
	.B1(N275),
	.A2(n494),
	.A1(n19), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U711 (
	.ZN(\regIn[12][15] ),
	.B2(n504),
	.B1(N275),
	.A2(n494),
	.A1(n21), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U712 (
	.ZN(\regIn[12][14] ),
	.B2(n505),
	.B1(N275),
	.A2(n494),
	.A1(n23), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U713 (
	.ZN(\regIn[12][13] ),
	.B2(n506),
	.B1(N275),
	.A2(n494),
	.A1(n25), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U714 (
	.ZN(\regIn[12][12] ),
	.B2(n507),
	.B1(N275),
	.A2(n494),
	.A1(n27), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U715 (
	.ZN(\regIn[12][11] ),
	.B2(n508),
	.B1(N275),
	.A2(n494),
	.A1(n29), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U716 (
	.ZN(\regIn[12][10] ),
	.B2(n509),
	.B1(N275),
	.A2(n494),
	.A1(n31), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U717 (
	.ZN(\regIn[12][0] ),
	.B2(n510),
	.B1(N275),
	.A2(n494),
	.A1(n33), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U718 (
	.ZN(n494),
	.A(N275), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U719 (
	.ZN(\regIn[11][9] ),
	.A(n511), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U720 (
	.ZN(n511),
	.B2(\regOut[11][9] ),
	.B1(n512),
	.A2(N269),
	.A1(dataIn[9]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U721 (
	.ZN(\regIn[11][8] ),
	.A(n513), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U722 (
	.ZN(n513),
	.B2(\regOut[11][8] ),
	.B1(n512),
	.A2(N269),
	.A1(dataIn[8]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U723 (
	.ZN(\regIn[11][7] ),
	.A(n514), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U724 (
	.ZN(n514),
	.B2(\regOut[11][7] ),
	.B1(n512),
	.A2(N269),
	.A1(dataIn[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U725 (
	.ZN(\regIn[11][6] ),
	.A(n515), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U726 (
	.ZN(n515),
	.B2(\regOut[11][6] ),
	.B1(n512),
	.A2(N269),
	.A1(dataIn[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U727 (
	.ZN(\regIn[11][5] ),
	.A(n516), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U728 (
	.ZN(n516),
	.B2(\regOut[11][5] ),
	.B1(n512),
	.A2(N269),
	.A1(dataIn[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U729 (
	.ZN(\regIn[11][4] ),
	.A(n517), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U730 (
	.ZN(n517),
	.B2(\regOut[11][4] ),
	.B1(n512),
	.A2(N269),
	.A1(dataIn[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U731 (
	.ZN(\regIn[11][3] ),
	.A(n518), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U732 (
	.ZN(n518),
	.B2(\regOut[11][3] ),
	.B1(n512),
	.A2(N269),
	.A1(dataIn[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U733 (
	.ZN(\regIn[11][2] ),
	.A(n519), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U734 (
	.ZN(n519),
	.B2(\regOut[11][2] ),
	.B1(n512),
	.A2(N269),
	.A1(dataIn[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U735 (
	.ZN(\regIn[11][1] ),
	.A(n520), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U736 (
	.ZN(n520),
	.B2(\regOut[11][1] ),
	.B1(n512),
	.A2(N269),
	.A1(dataIn[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U737 (
	.ZN(\regIn[11][15] ),
	.A(n521), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U738 (
	.ZN(n521),
	.B2(\regOut[11][15] ),
	.B1(n512),
	.A2(N269),
	.A1(dataIn[15]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U739 (
	.ZN(\regIn[11][14] ),
	.A(n522), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U740 (
	.ZN(n522),
	.B2(\regOut[11][14] ),
	.B1(n512),
	.A2(N269),
	.A1(dataIn[14]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U741 (
	.ZN(\regIn[11][13] ),
	.A(n523), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U742 (
	.ZN(n523),
	.B2(\regOut[11][13] ),
	.B1(n512),
	.A2(N269),
	.A1(dataIn[13]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U743 (
	.ZN(\regIn[11][12] ),
	.A(n524), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U744 (
	.ZN(n524),
	.B2(\regOut[11][12] ),
	.B1(n512),
	.A2(N269),
	.A1(dataIn[12]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U745 (
	.ZN(\regIn[11][11] ),
	.A(n525), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U746 (
	.ZN(n525),
	.B2(\regOut[11][11] ),
	.B1(n512),
	.A2(N269),
	.A1(dataIn[11]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U747 (
	.ZN(\regIn[11][10] ),
	.A(n526), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U748 (
	.ZN(n526),
	.B2(\regOut[11][10] ),
	.B1(n512),
	.A2(N269),
	.A1(dataIn[10]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U749 (
	.ZN(\regIn[11][0] ),
	.A(n527), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U750 (
	.ZN(n527),
	.B2(\regOut[11][0] ),
	.B1(n512),
	.A2(N269),
	.A1(dataIn[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U751 (
	.ZN(n512),
	.A(N269), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U752 (
	.ZN(\regIn[10][9] ),
	.A(n528), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U753 (
	.ZN(n528),
	.B2(\regOut[10][9] ),
	.B1(n529),
	.A2(N263),
	.A1(dataIn[9]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U754 (
	.ZN(\regIn[10][8] ),
	.A(n530), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U755 (
	.ZN(n530),
	.B2(\regOut[10][8] ),
	.B1(n529),
	.A2(N263),
	.A1(dataIn[8]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U756 (
	.ZN(\regIn[10][7] ),
	.A(n531), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U757 (
	.ZN(n531),
	.B2(\regOut[10][7] ),
	.B1(n529),
	.A2(N263),
	.A1(dataIn[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U758 (
	.ZN(\regIn[10][6] ),
	.A(n532), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U759 (
	.ZN(n532),
	.B2(\regOut[10][6] ),
	.B1(n529),
	.A2(N263),
	.A1(dataIn[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U760 (
	.ZN(\regIn[10][5] ),
	.A(n533), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U761 (
	.ZN(n533),
	.B2(\regOut[10][5] ),
	.B1(n529),
	.A2(N263),
	.A1(dataIn[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U762 (
	.ZN(\regIn[10][4] ),
	.A(n534), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U763 (
	.ZN(n534),
	.B2(\regOut[10][4] ),
	.B1(n529),
	.A2(N263),
	.A1(dataIn[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U764 (
	.ZN(\regIn[10][3] ),
	.A(n535), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U765 (
	.ZN(n535),
	.B2(\regOut[10][3] ),
	.B1(n529),
	.A2(N263),
	.A1(dataIn[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U766 (
	.ZN(\regIn[10][2] ),
	.A(n536), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U767 (
	.ZN(n536),
	.B2(\regOut[10][2] ),
	.B1(n529),
	.A2(N263),
	.A1(dataIn[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U768 (
	.ZN(\regIn[10][1] ),
	.A(n537), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U769 (
	.ZN(n537),
	.B2(\regOut[10][1] ),
	.B1(n529),
	.A2(N263),
	.A1(dataIn[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U770 (
	.ZN(\regIn[10][15] ),
	.A(n538), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U771 (
	.ZN(n538),
	.B2(\regOut[10][15] ),
	.B1(n529),
	.A2(N263),
	.A1(dataIn[15]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U772 (
	.ZN(\regIn[10][14] ),
	.A(n539), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U773 (
	.ZN(n539),
	.B2(\regOut[10][14] ),
	.B1(n529),
	.A2(N263),
	.A1(dataIn[14]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U774 (
	.ZN(\regIn[10][13] ),
	.A(n540), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U775 (
	.ZN(n540),
	.B2(\regOut[10][13] ),
	.B1(n529),
	.A2(N263),
	.A1(dataIn[13]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U776 (
	.ZN(\regIn[10][12] ),
	.A(n541), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U777 (
	.ZN(n541),
	.B2(\regOut[10][12] ),
	.B1(n529),
	.A2(N263),
	.A1(dataIn[12]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U778 (
	.ZN(\regIn[10][11] ),
	.A(n542), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U779 (
	.ZN(n542),
	.B2(\regOut[10][11] ),
	.B1(n529),
	.A2(N263),
	.A1(dataIn[11]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U780 (
	.ZN(\regIn[10][10] ),
	.A(n543), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U781 (
	.ZN(n543),
	.B2(\regOut[10][10] ),
	.B1(n529),
	.A2(N263),
	.A1(dataIn[10]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U782 (
	.ZN(\regIn[10][0] ),
	.A(n544), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U783 (
	.ZN(n544),
	.B2(\regOut[10][0] ),
	.B1(n529),
	.A2(N263),
	.A1(dataIn[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U784 (
	.ZN(n529),
	.A(N263), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U785 (
	.ZN(\regIn[0][9] ),
	.B2(n546),
	.B1(N199),
	.A2(n545),
	.A1(n3), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X2 U786 (
	.ZN(n3),
	.A(dataIn[9]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U787 (
	.ZN(\regIn[0][8] ),
	.B2(n547),
	.B1(N199),
	.A2(n545),
	.A1(n5), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X2 U788 (
	.ZN(n5),
	.A(dataIn[8]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U789 (
	.ZN(\regIn[0][7] ),
	.B2(n548),
	.B1(N199),
	.A2(n545),
	.A1(n7), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X2 U790 (
	.ZN(n7),
	.A(dataIn[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U791 (
	.ZN(\regIn[0][6] ),
	.B2(n549),
	.B1(N199),
	.A2(n545),
	.A1(n9), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X2 U792 (
	.ZN(n9),
	.A(dataIn[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U793 (
	.ZN(\regIn[0][5] ),
	.B2(n550),
	.B1(N199),
	.A2(n545),
	.A1(n11), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X2 U794 (
	.ZN(n11),
	.A(dataIn[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U795 (
	.ZN(\regIn[0][4] ),
	.B2(n551),
	.B1(N199),
	.A2(n545),
	.A1(n13), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X2 U796 (
	.ZN(n13),
	.A(dataIn[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U797 (
	.ZN(\regIn[0][3] ),
	.B2(n552),
	.B1(N199),
	.A2(n545),
	.A1(n15), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X2 U798 (
	.ZN(n15),
	.A(dataIn[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U799 (
	.ZN(\regIn[0][2] ),
	.B2(n553),
	.B1(N199),
	.A2(n545),
	.A1(n17), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X2 U800 (
	.ZN(n17),
	.A(dataIn[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U801 (
	.ZN(\regIn[0][1] ),
	.B2(n554),
	.B1(N199),
	.A2(n545),
	.A1(n19), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X2 U802 (
	.ZN(n19),
	.A(dataIn[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U803 (
	.ZN(\regIn[0][15] ),
	.B2(n555),
	.B1(N199),
	.A2(n545),
	.A1(n21), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X2 U804 (
	.ZN(n21),
	.A(dataIn[15]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U805 (
	.ZN(\regIn[0][14] ),
	.B2(n556),
	.B1(N199),
	.A2(n545),
	.A1(n23), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X2 U806 (
	.ZN(n23),
	.A(dataIn[14]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U807 (
	.ZN(\regIn[0][13] ),
	.B2(n557),
	.B1(N199),
	.A2(n545),
	.A1(n25), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X2 U808 (
	.ZN(n25),
	.A(dataIn[13]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U809 (
	.ZN(\regIn[0][12] ),
	.B2(n558),
	.B1(N199),
	.A2(n545),
	.A1(n27), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X2 U810 (
	.ZN(n27),
	.A(dataIn[12]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U811 (
	.ZN(\regIn[0][11] ),
	.B2(n559),
	.B1(N199),
	.A2(n545),
	.A1(n29), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X2 U812 (
	.ZN(n29),
	.A(dataIn[11]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U813 (
	.ZN(\regIn[0][10] ),
	.B2(n560),
	.B1(N199),
	.A2(n545),
	.A1(n31), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X2 U814 (
	.ZN(n31),
	.A(dataIn[10]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22_X1 U815 (
	.ZN(\regIn[0][0] ),
	.B2(n561),
	.B1(N199),
	.A2(n545),
	.A1(n33), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U816 (
	.ZN(n545),
	.A(N199), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X2 U817 (
	.ZN(n33),
	.A(dataIn[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U818 (
	.ZN(outB[9]),
	.A2(n563),
	.A1(n562), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4_X1 U819 (
	.ZN(n563),
	.A4(n567),
	.A3(n566),
	.A2(n565),
	.A1(n564), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U820 (
	.ZN(n567),
	.C2(FE_OFN75_n569),
	.C1(n427),
	.B2(FE_OFN74_n568),
	.B1(n410),
	.A(n570), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U821 (
	.ZN(n570),
	.B2(\regOut[18][9] ),
	.B1(n572),
	.A2(\regOut[19][9] ),
	.A1(n571), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U822 (
	.ZN(n566),
	.C2(FE_OFN73_n574),
	.C1(n342),
	.B2(FE_OFN72_n573),
	.B1(n325),
	.A(n575), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U823 (
	.ZN(n575),
	.B2(\regOut[22][9] ),
	.B1(n577),
	.A2(\regOut[23][9] ),
	.A1(n576), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U824 (
	.ZN(n565),
	.C2(FE_OFN67_n579),
	.C1(n274),
	.B2(FE_OFN66_n578),
	.B1(n257),
	.A(n580), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U825 (
	.ZN(n580),
	.B2(\regOut[26][9] ),
	.B1(n582),
	.A2(\regOut[27][9] ),
	.A1(n581), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U826 (
	.ZN(n564),
	.C2(FE_OFN65_n584),
	.C1(n155),
	.B2(FE_OFN64_n583),
	.B1(n138),
	.A(n585), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U827 (
	.ZN(n585),
	.B2(\regOut[28][9] ),
	.B1(n587),
	.A2(\regOut[29][9] ),
	.A1(n586), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4_X1 U828 (
	.ZN(n562),
	.A4(n591),
	.A3(n590),
	.A2(n589),
	.A1(n588), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U829 (
	.ZN(n591),
	.C2(FE_OFN63_n593),
	.C1(n546),
	.B2(FE_OFN62_n592),
	.B1(n359),
	.A(n594), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U830 (
	.ZN(n594),
	.B2(\regOut[2][9] ),
	.B1(n596),
	.A2(\regOut[3][9] ),
	.A1(n595), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U831 (
	.ZN(n590),
	.C2(FE_OFN61_n598),
	.C1(n104),
	.B2(FE_OFN60_n597),
	.B1(n87),
	.A(n599), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U832 (
	.ZN(n599),
	.B2(\regOut[6][9] ),
	.B1(n601),
	.A2(\regOut[7][9] ),
	.A1(n600), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U833 (
	.ZN(n589),
	.C2(FE_OFN71_n603),
	.C1(n36),
	.B2(FE_OFN70_n602),
	.B1(n4),
	.A(n604), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U834 (
	.ZN(n604),
	.B2(\regOut[10][9] ),
	.B1(n606),
	.A2(\regOut[11][9] ),
	.A1(n605), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U835 (
	.ZN(n588),
	.C2(FE_OFN69_n608),
	.C1(n495),
	.B2(FE_OFN68_n607),
	.B1(n478),
	.A(n609), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U836 (
	.ZN(n609),
	.B2(\regOut[14][9] ),
	.B1(n611),
	.A2(\regOut[15][9] ),
	.A1(n610), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U837 (
	.ZN(outB[8]),
	.A2(n613),
	.A1(n612), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4_X1 U838 (
	.ZN(n613),
	.A4(n617),
	.A3(n616),
	.A2(n615),
	.A1(n614), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U839 (
	.ZN(n617),
	.C2(FE_OFN75_n569),
	.C1(n428),
	.B2(FE_OFN74_n568),
	.B1(n411),
	.A(n618), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U840 (
	.ZN(n618),
	.B2(\regOut[18][8] ),
	.B1(n572),
	.A2(\regOut[19][8] ),
	.A1(n571), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U841 (
	.ZN(n616),
	.C2(FE_OFN73_n574),
	.C1(n343),
	.B2(FE_OFN72_n573),
	.B1(n326),
	.A(n619), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U842 (
	.ZN(n619),
	.B2(\regOut[22][8] ),
	.B1(n577),
	.A2(\regOut[23][8] ),
	.A1(n576), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U843 (
	.ZN(n615),
	.C2(FE_OFN67_n579),
	.C1(n275),
	.B2(FE_OFN66_n578),
	.B1(n258),
	.A(n620), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U844 (
	.ZN(n620),
	.B2(\regOut[26][8] ),
	.B1(n582),
	.A2(\regOut[27][8] ),
	.A1(n581), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U845 (
	.ZN(n614),
	.C2(FE_OFN65_n584),
	.C1(n156),
	.B2(FE_OFN64_n583),
	.B1(n139),
	.A(n621), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U846 (
	.ZN(n621),
	.B2(\regOut[28][8] ),
	.B1(n587),
	.A2(\regOut[29][8] ),
	.A1(n586), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4_X1 U847 (
	.ZN(n612),
	.A4(n625),
	.A3(n624),
	.A2(n623),
	.A1(n622), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U848 (
	.ZN(n625),
	.C2(FE_OFN63_n593),
	.C1(n547),
	.B2(FE_OFN62_n592),
	.B1(n360),
	.A(n626), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U849 (
	.ZN(n626),
	.B2(\regOut[2][8] ),
	.B1(n596),
	.A2(\regOut[3][8] ),
	.A1(n595), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U850 (
	.ZN(n624),
	.C2(FE_OFN61_n598),
	.C1(n105),
	.B2(FE_OFN60_n597),
	.B1(n88),
	.A(n627), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U851 (
	.ZN(n627),
	.B2(\regOut[6][8] ),
	.B1(n601),
	.A2(\regOut[7][8] ),
	.A1(n600), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U852 (
	.ZN(n623),
	.C2(FE_OFN71_n603),
	.C1(n37),
	.B2(FE_OFN70_n602),
	.B1(n6),
	.A(n628), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U853 (
	.ZN(n628),
	.B2(\regOut[10][8] ),
	.B1(n606),
	.A2(\regOut[11][8] ),
	.A1(n605), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U854 (
	.ZN(n622),
	.C2(FE_OFN69_n608),
	.C1(n496),
	.B2(FE_OFN68_n607),
	.B1(n479),
	.A(n629), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U855 (
	.ZN(n629),
	.B2(\regOut[14][8] ),
	.B1(n611),
	.A2(\regOut[15][8] ),
	.A1(n610), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U856 (
	.ZN(outB[7]),
	.A2(n631),
	.A1(n630), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4_X1 U857 (
	.ZN(n631),
	.A4(n635),
	.A3(n634),
	.A2(n633),
	.A1(n632), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U858 (
	.ZN(n635),
	.C2(FE_OFN75_n569),
	.C1(n429),
	.B2(FE_OFN74_n568),
	.B1(n412),
	.A(n636), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U859 (
	.ZN(n636),
	.B2(\regOut[18][7] ),
	.B1(n572),
	.A2(\regOut[19][7] ),
	.A1(n571), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U860 (
	.ZN(n634),
	.C2(FE_OFN73_n574),
	.C1(n344),
	.B2(FE_OFN72_n573),
	.B1(n327),
	.A(n637), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U861 (
	.ZN(n637),
	.B2(\regOut[22][7] ),
	.B1(n577),
	.A2(\regOut[23][7] ),
	.A1(n576), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U862 (
	.ZN(n633),
	.C2(FE_OFN67_n579),
	.C1(n276),
	.B2(FE_OFN66_n578),
	.B1(n259),
	.A(n638), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U863 (
	.ZN(n638),
	.B2(\regOut[26][7] ),
	.B1(n582),
	.A2(\regOut[27][7] ),
	.A1(n581), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U864 (
	.ZN(n632),
	.C2(FE_OFN65_n584),
	.C1(n157),
	.B2(FE_OFN64_n583),
	.B1(n140),
	.A(n639), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U865 (
	.ZN(n639),
	.B2(\regOut[28][7] ),
	.B1(n587),
	.A2(\regOut[29][7] ),
	.A1(n586), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4_X1 U866 (
	.ZN(n630),
	.A4(n643),
	.A3(n642),
	.A2(n641),
	.A1(n640), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U867 (
	.ZN(n643),
	.C2(FE_OFN63_n593),
	.C1(n548),
	.B2(FE_OFN62_n592),
	.B1(n361),
	.A(n644), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U868 (
	.ZN(n644),
	.B2(\regOut[2][7] ),
	.B1(n596),
	.A2(\regOut[3][7] ),
	.A1(n595), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U869 (
	.ZN(n642),
	.C2(FE_OFN61_n598),
	.C1(n106),
	.B2(FE_OFN60_n597),
	.B1(n89),
	.A(n645), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U870 (
	.ZN(n645),
	.B2(\regOut[6][7] ),
	.B1(n601),
	.A2(\regOut[7][7] ),
	.A1(n600), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U871 (
	.ZN(n641),
	.C2(FE_OFN71_n603),
	.C1(n38),
	.B2(FE_OFN70_n602),
	.B1(n8),
	.A(n646), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U872 (
	.ZN(n646),
	.B2(\regOut[10][7] ),
	.B1(n606),
	.A2(\regOut[11][7] ),
	.A1(n605), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U873 (
	.ZN(n640),
	.C2(FE_OFN69_n608),
	.C1(n497),
	.B2(FE_OFN68_n607),
	.B1(n480),
	.A(n647), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U874 (
	.ZN(n647),
	.B2(\regOut[14][7] ),
	.B1(n611),
	.A2(\regOut[15][7] ),
	.A1(n610), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U875 (
	.ZN(outB[6]),
	.A2(n649),
	.A1(n648), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4_X1 U876 (
	.ZN(n649),
	.A4(n653),
	.A3(n652),
	.A2(n651),
	.A1(n650), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U877 (
	.ZN(n653),
	.C2(FE_OFN75_n569),
	.C1(n430),
	.B2(FE_OFN74_n568),
	.B1(n413),
	.A(n654), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U878 (
	.ZN(n654),
	.B2(\regOut[18][6] ),
	.B1(n572),
	.A2(\regOut[19][6] ),
	.A1(n571), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U879 (
	.ZN(n652),
	.C2(FE_OFN73_n574),
	.C1(n345),
	.B2(FE_OFN72_n573),
	.B1(n328),
	.A(n655), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U880 (
	.ZN(n655),
	.B2(\regOut[22][6] ),
	.B1(n577),
	.A2(\regOut[23][6] ),
	.A1(n576), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U881 (
	.ZN(n651),
	.C2(FE_OFN67_n579),
	.C1(n277),
	.B2(FE_OFN66_n578),
	.B1(n260),
	.A(n656), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U882 (
	.ZN(n656),
	.B2(\regOut[26][6] ),
	.B1(n582),
	.A2(\regOut[27][6] ),
	.A1(n581), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U883 (
	.ZN(n650),
	.C2(FE_OFN65_n584),
	.C1(n158),
	.B2(FE_OFN64_n583),
	.B1(n141),
	.A(n657), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U884 (
	.ZN(n657),
	.B2(\regOut[28][6] ),
	.B1(n587),
	.A2(\regOut[29][6] ),
	.A1(n586), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4_X1 U885 (
	.ZN(n648),
	.A4(n661),
	.A3(n660),
	.A2(n659),
	.A1(n658), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U886 (
	.ZN(n661),
	.C2(FE_OFN63_n593),
	.C1(n549),
	.B2(FE_OFN62_n592),
	.B1(n362),
	.A(n662), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U887 (
	.ZN(n662),
	.B2(\regOut[2][6] ),
	.B1(n596),
	.A2(\regOut[3][6] ),
	.A1(n595), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U888 (
	.ZN(n660),
	.C2(FE_OFN61_n598),
	.C1(n107),
	.B2(FE_OFN60_n597),
	.B1(n90),
	.A(n663), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U889 (
	.ZN(n663),
	.B2(\regOut[6][6] ),
	.B1(n601),
	.A2(\regOut[7][6] ),
	.A1(n600), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U890 (
	.ZN(n659),
	.C2(FE_OFN71_n603),
	.C1(n39),
	.B2(FE_OFN70_n602),
	.B1(n10),
	.A(n664), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U891 (
	.ZN(n664),
	.B2(\regOut[10][6] ),
	.B1(n606),
	.A2(\regOut[11][6] ),
	.A1(n605), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U892 (
	.ZN(n658),
	.C2(FE_OFN69_n608),
	.C1(n498),
	.B2(FE_OFN68_n607),
	.B1(n481),
	.A(n665), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U893 (
	.ZN(n665),
	.B2(\regOut[14][6] ),
	.B1(n611),
	.A2(\regOut[15][6] ),
	.A1(n610), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U894 (
	.ZN(outB[5]),
	.A2(n667),
	.A1(n666), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4_X1 U895 (
	.ZN(n667),
	.A4(n671),
	.A3(n670),
	.A2(n669),
	.A1(n668), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U896 (
	.ZN(n671),
	.C2(FE_OFN75_n569),
	.C1(n431),
	.B2(FE_OFN74_n568),
	.B1(n414),
	.A(n672), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U897 (
	.ZN(n672),
	.B2(\regOut[18][5] ),
	.B1(n572),
	.A2(\regOut[19][5] ),
	.A1(n571), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U898 (
	.ZN(n670),
	.C2(FE_OFN73_n574),
	.C1(n346),
	.B2(FE_OFN72_n573),
	.B1(n329),
	.A(n673), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U899 (
	.ZN(n673),
	.B2(\regOut[22][5] ),
	.B1(n577),
	.A2(\regOut[23][5] ),
	.A1(n576), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U900 (
	.ZN(n669),
	.C2(FE_OFN67_n579),
	.C1(n278),
	.B2(FE_OFN66_n578),
	.B1(n261),
	.A(n674), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U901 (
	.ZN(n674),
	.B2(\regOut[26][5] ),
	.B1(n582),
	.A2(\regOut[27][5] ),
	.A1(n581), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U902 (
	.ZN(n668),
	.C2(FE_OFN65_n584),
	.C1(n159),
	.B2(FE_OFN64_n583),
	.B1(n142),
	.A(n675), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U903 (
	.ZN(n675),
	.B2(\regOut[28][5] ),
	.B1(n587),
	.A2(\regOut[29][5] ),
	.A1(n586), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4_X1 U904 (
	.ZN(n666),
	.A4(n679),
	.A3(n678),
	.A2(n677),
	.A1(n676), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U905 (
	.ZN(n679),
	.C2(FE_OFN63_n593),
	.C1(n550),
	.B2(FE_OFN62_n592),
	.B1(n363),
	.A(n680), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U906 (
	.ZN(n680),
	.B2(\regOut[2][5] ),
	.B1(n596),
	.A2(\regOut[3][5] ),
	.A1(n595), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U907 (
	.ZN(n678),
	.C2(FE_OFN61_n598),
	.C1(n108),
	.B2(FE_OFN60_n597),
	.B1(n91),
	.A(n681), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U908 (
	.ZN(n681),
	.B2(\regOut[6][5] ),
	.B1(n601),
	.A2(\regOut[7][5] ),
	.A1(n600), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U909 (
	.ZN(n677),
	.C2(FE_OFN71_n603),
	.C1(n40),
	.B2(FE_OFN70_n602),
	.B1(n12),
	.A(n682), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U910 (
	.ZN(n682),
	.B2(\regOut[10][5] ),
	.B1(n606),
	.A2(\regOut[11][5] ),
	.A1(n605), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U911 (
	.ZN(n676),
	.C2(FE_OFN69_n608),
	.C1(n499),
	.B2(FE_OFN68_n607),
	.B1(n482),
	.A(n683), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U912 (
	.ZN(n683),
	.B2(\regOut[14][5] ),
	.B1(n611),
	.A2(\regOut[15][5] ),
	.A1(n610), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U913 (
	.ZN(outB[4]),
	.A2(n685),
	.A1(n684), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4_X1 U914 (
	.ZN(n685),
	.A4(n689),
	.A3(n688),
	.A2(n687),
	.A1(n686), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U915 (
	.ZN(n689),
	.C2(FE_OFN75_n569),
	.C1(n432),
	.B2(FE_OFN74_n568),
	.B1(n415),
	.A(n690), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U916 (
	.ZN(n690),
	.B2(\regOut[18][4] ),
	.B1(n572),
	.A2(\regOut[19][4] ),
	.A1(n571), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U917 (
	.ZN(n688),
	.C2(FE_OFN73_n574),
	.C1(n347),
	.B2(FE_OFN72_n573),
	.B1(n330),
	.A(n691), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U918 (
	.ZN(n691),
	.B2(\regOut[22][4] ),
	.B1(n577),
	.A2(\regOut[23][4] ),
	.A1(n576), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U919 (
	.ZN(n687),
	.C2(FE_OFN67_n579),
	.C1(n279),
	.B2(FE_OFN66_n578),
	.B1(n262),
	.A(n692), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U920 (
	.ZN(n692),
	.B2(\regOut[26][4] ),
	.B1(n582),
	.A2(\regOut[27][4] ),
	.A1(n581), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U921 (
	.ZN(n686),
	.C2(FE_OFN65_n584),
	.C1(n160),
	.B2(FE_OFN64_n583),
	.B1(n143),
	.A(n693), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U922 (
	.ZN(n693),
	.B2(\regOut[28][4] ),
	.B1(n587),
	.A2(\regOut[29][4] ),
	.A1(n586), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4_X1 U923 (
	.ZN(n684),
	.A4(n697),
	.A3(n696),
	.A2(n695),
	.A1(n694), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U924 (
	.ZN(n697),
	.C2(FE_OFN63_n593),
	.C1(n551),
	.B2(FE_OFN62_n592),
	.B1(n364),
	.A(n698), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U925 (
	.ZN(n698),
	.B2(\regOut[2][4] ),
	.B1(n596),
	.A2(\regOut[3][4] ),
	.A1(n595), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U926 (
	.ZN(n696),
	.C2(FE_OFN61_n598),
	.C1(n109),
	.B2(FE_OFN60_n597),
	.B1(n92),
	.A(n699), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U927 (
	.ZN(n699),
	.B2(\regOut[6][4] ),
	.B1(n601),
	.A2(\regOut[7][4] ),
	.A1(n600), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U928 (
	.ZN(n695),
	.C2(FE_OFN71_n603),
	.C1(n41),
	.B2(FE_OFN70_n602),
	.B1(n14),
	.A(n700), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U929 (
	.ZN(n700),
	.B2(\regOut[10][4] ),
	.B1(n606),
	.A2(\regOut[11][4] ),
	.A1(n605), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U930 (
	.ZN(n694),
	.C2(FE_OFN69_n608),
	.C1(n500),
	.B2(FE_OFN68_n607),
	.B1(n483),
	.A(n701), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U931 (
	.ZN(n701),
	.B2(\regOut[14][4] ),
	.B1(n611),
	.A2(\regOut[15][4] ),
	.A1(n610), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U932 (
	.ZN(outB[3]),
	.A2(n703),
	.A1(n702), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4_X1 U933 (
	.ZN(n703),
	.A4(n707),
	.A3(n706),
	.A2(n705),
	.A1(n704), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U934 (
	.ZN(n707),
	.C2(FE_OFN75_n569),
	.C1(n433),
	.B2(FE_OFN74_n568),
	.B1(n416),
	.A(n708), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U935 (
	.ZN(n708),
	.B2(\regOut[18][3] ),
	.B1(n572),
	.A2(\regOut[19][3] ),
	.A1(n571), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U936 (
	.ZN(n706),
	.C2(FE_OFN73_n574),
	.C1(n348),
	.B2(FE_OFN72_n573),
	.B1(n331),
	.A(n709), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U937 (
	.ZN(n709),
	.B2(\regOut[22][3] ),
	.B1(n577),
	.A2(\regOut[23][3] ),
	.A1(n576), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U938 (
	.ZN(n705),
	.C2(FE_OFN67_n579),
	.C1(n280),
	.B2(FE_OFN66_n578),
	.B1(n263),
	.A(n710), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U939 (
	.ZN(n710),
	.B2(\regOut[26][3] ),
	.B1(n582),
	.A2(\regOut[27][3] ),
	.A1(n581), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U940 (
	.ZN(n704),
	.C2(FE_OFN65_n584),
	.C1(n161),
	.B2(FE_OFN64_n583),
	.B1(n144),
	.A(n711), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U941 (
	.ZN(n711),
	.B2(\regOut[28][3] ),
	.B1(n587),
	.A2(\regOut[29][3] ),
	.A1(n586), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4_X1 U942 (
	.ZN(n702),
	.A4(n715),
	.A3(n714),
	.A2(n713),
	.A1(n712), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U943 (
	.ZN(n715),
	.C2(FE_OFN63_n593),
	.C1(n552),
	.B2(FE_OFN62_n592),
	.B1(n365),
	.A(n716), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U944 (
	.ZN(n716),
	.B2(\regOut[2][3] ),
	.B1(n596),
	.A2(\regOut[3][3] ),
	.A1(n595), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U945 (
	.ZN(n714),
	.C2(FE_OFN61_n598),
	.C1(n110),
	.B2(FE_OFN60_n597),
	.B1(n93),
	.A(n717), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U946 (
	.ZN(n717),
	.B2(\regOut[6][3] ),
	.B1(n601),
	.A2(\regOut[7][3] ),
	.A1(n600), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U947 (
	.ZN(n713),
	.C2(FE_OFN71_n603),
	.C1(n42),
	.B2(n602),
	.B1(n16),
	.A(n718), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U948 (
	.ZN(n718),
	.B2(\regOut[10][3] ),
	.B1(n606),
	.A2(\regOut[11][3] ),
	.A1(n605), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U949 (
	.ZN(n712),
	.C2(FE_OFN69_n608),
	.C1(n501),
	.B2(FE_OFN68_n607),
	.B1(n484),
	.A(n719), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U950 (
	.ZN(n719),
	.B2(\regOut[14][3] ),
	.B1(n611),
	.A2(\regOut[15][3] ),
	.A1(n610), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U951 (
	.ZN(outB[2]),
	.A2(n721),
	.A1(n720), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4_X1 U952 (
	.ZN(n721),
	.A4(n725),
	.A3(n724),
	.A2(n723),
	.A1(n722), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U953 (
	.ZN(n725),
	.C2(FE_OFN75_n569),
	.C1(n434),
	.B2(FE_OFN74_n568),
	.B1(n417),
	.A(n726), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U954 (
	.ZN(n726),
	.B2(\regOut[18][2] ),
	.B1(n572),
	.A2(\regOut[19][2] ),
	.A1(n571), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U955 (
	.ZN(n724),
	.C2(FE_OFN73_n574),
	.C1(n349),
	.B2(FE_OFN72_n573),
	.B1(n332),
	.A(n727), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U956 (
	.ZN(n727),
	.B2(\regOut[22][2] ),
	.B1(n577),
	.A2(\regOut[23][2] ),
	.A1(n576), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U957 (
	.ZN(n723),
	.C2(FE_OFN67_n579),
	.C1(n281),
	.B2(FE_OFN66_n578),
	.B1(n264),
	.A(n728), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U958 (
	.ZN(n728),
	.B2(\regOut[26][2] ),
	.B1(n582),
	.A2(\regOut[27][2] ),
	.A1(n581), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U959 (
	.ZN(n722),
	.C2(FE_OFN65_n584),
	.C1(n162),
	.B2(FE_OFN64_n583),
	.B1(n145),
	.A(n729), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U960 (
	.ZN(n729),
	.B2(\regOut[28][2] ),
	.B1(n587),
	.A2(\regOut[29][2] ),
	.A1(n586), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4_X1 U961 (
	.ZN(n720),
	.A4(n733),
	.A3(n732),
	.A2(n731),
	.A1(n730), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U962 (
	.ZN(n733),
	.C2(FE_OFN63_n593),
	.C1(n553),
	.B2(FE_OFN62_n592),
	.B1(n366),
	.A(n734), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U963 (
	.ZN(n734),
	.B2(\regOut[2][2] ),
	.B1(n596),
	.A2(\regOut[3][2] ),
	.A1(n595), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U964 (
	.ZN(n732),
	.C2(FE_OFN61_n598),
	.C1(n111),
	.B2(FE_OFN60_n597),
	.B1(n94),
	.A(n735), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U965 (
	.ZN(n735),
	.B2(\regOut[6][2] ),
	.B1(n601),
	.A2(\regOut[7][2] ),
	.A1(n600), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U966 (
	.ZN(n731),
	.C2(FE_OFN71_n603),
	.C1(n43),
	.B2(FE_OFN70_n602),
	.B1(n18),
	.A(n736), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U967 (
	.ZN(n736),
	.B2(\regOut[10][2] ),
	.B1(n606),
	.A2(\regOut[11][2] ),
	.A1(n605), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U968 (
	.ZN(n730),
	.C2(FE_OFN69_n608),
	.C1(n502),
	.B2(FE_OFN68_n607),
	.B1(n485),
	.A(n737), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U969 (
	.ZN(n737),
	.B2(\regOut[14][2] ),
	.B1(n611),
	.A2(\regOut[15][2] ),
	.A1(n610), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U970 (
	.ZN(outB[1]),
	.A2(n739),
	.A1(n738), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4_X1 U971 (
	.ZN(n739),
	.A4(n743),
	.A3(n742),
	.A2(n741),
	.A1(n740), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U972 (
	.ZN(n743),
	.C2(FE_OFN75_n569),
	.C1(n435),
	.B2(FE_OFN74_n568),
	.B1(n418),
	.A(n744), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U973 (
	.ZN(n744),
	.B2(\regOut[18][1] ),
	.B1(n572),
	.A2(\regOut[19][1] ),
	.A1(n571), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U974 (
	.ZN(n742),
	.C2(FE_OFN73_n574),
	.C1(n350),
	.B2(FE_OFN72_n573),
	.B1(n333),
	.A(n745), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U975 (
	.ZN(n745),
	.B2(\regOut[22][1] ),
	.B1(n577),
	.A2(\regOut[23][1] ),
	.A1(n576), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U976 (
	.ZN(n741),
	.C2(FE_OFN67_n579),
	.C1(n282),
	.B2(FE_OFN66_n578),
	.B1(n265),
	.A(n746), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U977 (
	.ZN(n746),
	.B2(\regOut[26][1] ),
	.B1(n582),
	.A2(\regOut[27][1] ),
	.A1(n581), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U978 (
	.ZN(n740),
	.C2(FE_OFN65_n584),
	.C1(n163),
	.B2(FE_OFN64_n583),
	.B1(n146),
	.A(n747), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U979 (
	.ZN(n747),
	.B2(\regOut[28][1] ),
	.B1(n587),
	.A2(\regOut[29][1] ),
	.A1(n586), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4_X1 U980 (
	.ZN(n738),
	.A4(n751),
	.A3(n750),
	.A2(n749),
	.A1(n748), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U981 (
	.ZN(n751),
	.C2(FE_OFN63_n593),
	.C1(n554),
	.B2(FE_OFN62_n592),
	.B1(n367),
	.A(n752), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U982 (
	.ZN(n752),
	.B2(\regOut[2][1] ),
	.B1(n596),
	.A2(\regOut[3][1] ),
	.A1(n595), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U983 (
	.ZN(n750),
	.C2(FE_OFN61_n598),
	.C1(n112),
	.B2(FE_OFN60_n597),
	.B1(n95),
	.A(n753), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U984 (
	.ZN(n753),
	.B2(\regOut[6][1] ),
	.B1(n601),
	.A2(\regOut[7][1] ),
	.A1(n600), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U985 (
	.ZN(n749),
	.C2(FE_OFN71_n603),
	.C1(n44),
	.B2(FE_OFN70_n602),
	.B1(n20),
	.A(n754), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U986 (
	.ZN(n754),
	.B2(\regOut[10][1] ),
	.B1(n606),
	.A2(\regOut[11][1] ),
	.A1(n605), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U987 (
	.ZN(n748),
	.C2(FE_OFN69_n608),
	.C1(n503),
	.B2(FE_OFN68_n607),
	.B1(n486),
	.A(n755), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U988 (
	.ZN(n755),
	.B2(\regOut[14][1] ),
	.B1(n611),
	.A2(\regOut[15][1] ),
	.A1(n610), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U989 (
	.ZN(outB[15]),
	.A2(n757),
	.A1(n756), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4_X1 U990 (
	.ZN(n757),
	.A4(n761),
	.A3(n760),
	.A2(n759),
	.A1(n758), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U991 (
	.ZN(n761),
	.C2(FE_OFN75_n569),
	.C1(n436),
	.B2(FE_OFN74_n568),
	.B1(n419),
	.A(n762), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U992 (
	.ZN(n762),
	.B2(\regOut[18][15] ),
	.B1(n572),
	.A2(\regOut[19][15] ),
	.A1(n571), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U993 (
	.ZN(n760),
	.C2(FE_OFN73_n574),
	.C1(n351),
	.B2(FE_OFN72_n573),
	.B1(n334),
	.A(n763), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U994 (
	.ZN(n763),
	.B2(\regOut[22][15] ),
	.B1(n577),
	.A2(\regOut[23][15] ),
	.A1(n576), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U995 (
	.ZN(n759),
	.C2(FE_OFN67_n579),
	.C1(n283),
	.B2(FE_OFN66_n578),
	.B1(n266),
	.A(n764), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U996 (
	.ZN(n764),
	.B2(\regOut[26][15] ),
	.B1(n582),
	.A2(\regOut[27][15] ),
	.A1(n581), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U997 (
	.ZN(n758),
	.C2(FE_OFN65_n584),
	.C1(n164),
	.B2(FE_OFN64_n583),
	.B1(n147),
	.A(n765), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U998 (
	.ZN(n765),
	.B2(\regOut[28][15] ),
	.B1(n587),
	.A2(\regOut[29][15] ),
	.A1(n586), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4_X1 U999 (
	.ZN(n756),
	.A4(n769),
	.A3(n768),
	.A2(n767),
	.A1(n766), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U1000 (
	.ZN(n769),
	.C2(FE_OFN63_n593),
	.C1(n555),
	.B2(FE_OFN62_n592),
	.B1(n368),
	.A(n770), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U1001 (
	.ZN(n770),
	.B2(\regOut[2][15] ),
	.B1(n596),
	.A2(\regOut[3][15] ),
	.A1(n595), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U1002 (
	.ZN(n768),
	.C2(FE_OFN61_n598),
	.C1(n113),
	.B2(FE_OFN60_n597),
	.B1(n96),
	.A(n771), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U1003 (
	.ZN(n771),
	.B2(\regOut[6][15] ),
	.B1(n601),
	.A2(\regOut[7][15] ),
	.A1(n600), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U1004 (
	.ZN(n767),
	.C2(FE_OFN71_n603),
	.C1(n45),
	.B2(FE_OFN70_n602),
	.B1(n22),
	.A(n772), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U1005 (
	.ZN(n772),
	.B2(\regOut[10][15] ),
	.B1(n606),
	.A2(\regOut[11][15] ),
	.A1(n605), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U1006 (
	.ZN(n766),
	.C2(FE_OFN69_n608),
	.C1(n504),
	.B2(FE_OFN68_n607),
	.B1(n487),
	.A(n773), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U1007 (
	.ZN(n773),
	.B2(\regOut[14][15] ),
	.B1(n611),
	.A2(\regOut[15][15] ),
	.A1(n610), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U1008 (
	.ZN(outB[14]),
	.A2(n775),
	.A1(n774), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4_X1 U1009 (
	.ZN(n775),
	.A4(n779),
	.A3(n778),
	.A2(n777),
	.A1(n776), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U1010 (
	.ZN(n779),
	.C2(FE_OFN75_n569),
	.C1(n437),
	.B2(FE_OFN74_n568),
	.B1(n420),
	.A(n780), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U1011 (
	.ZN(n780),
	.B2(\regOut[18][14] ),
	.B1(n572),
	.A2(\regOut[19][14] ),
	.A1(n571), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U1012 (
	.ZN(n778),
	.C2(FE_OFN73_n574),
	.C1(n352),
	.B2(FE_OFN72_n573),
	.B1(n335),
	.A(n781), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U1013 (
	.ZN(n781),
	.B2(\regOut[22][14] ),
	.B1(n577),
	.A2(\regOut[23][14] ),
	.A1(n576), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U1014 (
	.ZN(n777),
	.C2(FE_OFN67_n579),
	.C1(n284),
	.B2(FE_OFN66_n578),
	.B1(n267),
	.A(n782), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U1015 (
	.ZN(n782),
	.B2(\regOut[26][14] ),
	.B1(n582),
	.A2(\regOut[27][14] ),
	.A1(n581), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U1016 (
	.ZN(n776),
	.C2(FE_OFN65_n584),
	.C1(n165),
	.B2(FE_OFN64_n583),
	.B1(n148),
	.A(n783), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U1017 (
	.ZN(n783),
	.B2(\regOut[28][14] ),
	.B1(n587),
	.A2(\regOut[29][14] ),
	.A1(n586), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4_X1 U1018 (
	.ZN(n774),
	.A4(n787),
	.A3(n786),
	.A2(n785),
	.A1(n784), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U1019 (
	.ZN(n787),
	.C2(FE_OFN63_n593),
	.C1(n556),
	.B2(FE_OFN62_n592),
	.B1(n369),
	.A(n788), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U1020 (
	.ZN(n788),
	.B2(\regOut[2][14] ),
	.B1(n596),
	.A2(\regOut[3][14] ),
	.A1(n595), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U1021 (
	.ZN(n786),
	.C2(FE_OFN61_n598),
	.C1(n114),
	.B2(FE_OFN60_n597),
	.B1(n97),
	.A(n789), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U1022 (
	.ZN(n789),
	.B2(\regOut[6][14] ),
	.B1(n601),
	.A2(\regOut[7][14] ),
	.A1(n600), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U1023 (
	.ZN(n785),
	.C2(FE_OFN71_n603),
	.C1(n46),
	.B2(FE_OFN70_n602),
	.B1(n24),
	.A(n790), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U1024 (
	.ZN(n790),
	.B2(\regOut[10][14] ),
	.B1(n606),
	.A2(\regOut[11][14] ),
	.A1(n605), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U1025 (
	.ZN(n784),
	.C2(FE_OFN69_n608),
	.C1(n505),
	.B2(FE_OFN68_n607),
	.B1(n488),
	.A(n791), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U1026 (
	.ZN(n791),
	.B2(\regOut[14][14] ),
	.B1(n611),
	.A2(\regOut[15][14] ),
	.A1(n610), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U1027 (
	.ZN(outB[13]),
	.A2(n793),
	.A1(n792), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4_X1 U1028 (
	.ZN(n793),
	.A4(n797),
	.A3(n796),
	.A2(n795),
	.A1(n794), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U1029 (
	.ZN(n797),
	.C2(FE_OFN75_n569),
	.C1(n438),
	.B2(FE_OFN74_n568),
	.B1(n421),
	.A(n798), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U1030 (
	.ZN(n798),
	.B2(\regOut[18][13] ),
	.B1(n572),
	.A2(\regOut[19][13] ),
	.A1(n571), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U1031 (
	.ZN(n796),
	.C2(FE_OFN73_n574),
	.C1(n353),
	.B2(FE_OFN72_n573),
	.B1(n336),
	.A(n799), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U1032 (
	.ZN(n799),
	.B2(\regOut[22][13] ),
	.B1(n577),
	.A2(\regOut[23][13] ),
	.A1(n576), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U1033 (
	.ZN(n795),
	.C2(FE_OFN67_n579),
	.C1(n285),
	.B2(FE_OFN66_n578),
	.B1(n268),
	.A(n800), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U1034 (
	.ZN(n800),
	.B2(\regOut[26][13] ),
	.B1(n582),
	.A2(\regOut[27][13] ),
	.A1(n581), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U1035 (
	.ZN(n794),
	.C2(FE_OFN65_n584),
	.C1(n166),
	.B2(FE_OFN64_n583),
	.B1(n149),
	.A(n801), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U1036 (
	.ZN(n801),
	.B2(\regOut[28][13] ),
	.B1(n587),
	.A2(\regOut[29][13] ),
	.A1(n586), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4_X1 U1037 (
	.ZN(n792),
	.A4(n805),
	.A3(n804),
	.A2(n803),
	.A1(n802), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U1038 (
	.ZN(n805),
	.C2(FE_OFN63_n593),
	.C1(n557),
	.B2(FE_OFN62_n592),
	.B1(n370),
	.A(n806), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U1039 (
	.ZN(n806),
	.B2(\regOut[2][13] ),
	.B1(n596),
	.A2(\regOut[3][13] ),
	.A1(n595), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U1040 (
	.ZN(n804),
	.C2(FE_OFN61_n598),
	.C1(n115),
	.B2(FE_OFN60_n597),
	.B1(n98),
	.A(n807), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U1041 (
	.ZN(n807),
	.B2(\regOut[6][13] ),
	.B1(n601),
	.A2(\regOut[7][13] ),
	.A1(n600), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U1042 (
	.ZN(n803),
	.C2(FE_OFN71_n603),
	.C1(n47),
	.B2(FE_OFN70_n602),
	.B1(n26),
	.A(n808), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U1043 (
	.ZN(n808),
	.B2(\regOut[10][13] ),
	.B1(n606),
	.A2(\regOut[11][13] ),
	.A1(n605), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U1044 (
	.ZN(n802),
	.C2(FE_OFN69_n608),
	.C1(n506),
	.B2(FE_OFN68_n607),
	.B1(n489),
	.A(n809), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U1045 (
	.ZN(n809),
	.B2(\regOut[14][13] ),
	.B1(n611),
	.A2(\regOut[15][13] ),
	.A1(n610), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U1046 (
	.ZN(outB[12]),
	.A2(n811),
	.A1(n810), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4_X1 U1047 (
	.ZN(n811),
	.A4(n815),
	.A3(n814),
	.A2(n813),
	.A1(n812), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U1048 (
	.ZN(n815),
	.C2(FE_OFN75_n569),
	.C1(n439),
	.B2(FE_OFN74_n568),
	.B1(n422),
	.A(n816), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U1049 (
	.ZN(n816),
	.B2(\regOut[18][12] ),
	.B1(n572),
	.A2(\regOut[19][12] ),
	.A1(n571), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U1050 (
	.ZN(n814),
	.C2(FE_OFN73_n574),
	.C1(n354),
	.B2(FE_OFN72_n573),
	.B1(n337),
	.A(n817), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U1051 (
	.ZN(n817),
	.B2(\regOut[22][12] ),
	.B1(n577),
	.A2(\regOut[23][12] ),
	.A1(n576), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U1052 (
	.ZN(n813),
	.C2(FE_OFN67_n579),
	.C1(n286),
	.B2(FE_OFN66_n578),
	.B1(n269),
	.A(n818), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U1053 (
	.ZN(n818),
	.B2(\regOut[26][12] ),
	.B1(n582),
	.A2(\regOut[27][12] ),
	.A1(n581), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U1054 (
	.ZN(n812),
	.C2(FE_OFN65_n584),
	.C1(n167),
	.B2(FE_OFN64_n583),
	.B1(n150),
	.A(n819), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U1055 (
	.ZN(n819),
	.B2(\regOut[28][12] ),
	.B1(n587),
	.A2(\regOut[29][12] ),
	.A1(n586), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4_X1 U1056 (
	.ZN(n810),
	.A4(n823),
	.A3(n822),
	.A2(n821),
	.A1(n820), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U1057 (
	.ZN(n823),
	.C2(FE_OFN63_n593),
	.C1(n558),
	.B2(FE_OFN62_n592),
	.B1(n371),
	.A(n824), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U1058 (
	.ZN(n824),
	.B2(\regOut[2][12] ),
	.B1(n596),
	.A2(\regOut[3][12] ),
	.A1(n595), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U1059 (
	.ZN(n822),
	.C2(FE_OFN61_n598),
	.C1(n116),
	.B2(FE_OFN60_n597),
	.B1(n99),
	.A(n825), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U1060 (
	.ZN(n825),
	.B2(\regOut[6][12] ),
	.B1(n601),
	.A2(\regOut[7][12] ),
	.A1(n600), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U1061 (
	.ZN(n821),
	.C2(FE_OFN71_n603),
	.C1(n48),
	.B2(FE_OFN70_n602),
	.B1(n28),
	.A(n826), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U1062 (
	.ZN(n826),
	.B2(\regOut[10][12] ),
	.B1(n606),
	.A2(\regOut[11][12] ),
	.A1(n605), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U1063 (
	.ZN(n820),
	.C2(FE_OFN69_n608),
	.C1(n507),
	.B2(FE_OFN68_n607),
	.B1(n490),
	.A(n827), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U1064 (
	.ZN(n827),
	.B2(\regOut[14][12] ),
	.B1(n611),
	.A2(\regOut[15][12] ),
	.A1(n610), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U1065 (
	.ZN(outB[11]),
	.A2(n829),
	.A1(n828), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4_X1 U1066 (
	.ZN(n829),
	.A4(n833),
	.A3(n832),
	.A2(n831),
	.A1(n830), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U1067 (
	.ZN(n833),
	.C2(FE_OFN75_n569),
	.C1(n440),
	.B2(FE_OFN74_n568),
	.B1(n423),
	.A(n834), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U1068 (
	.ZN(n834),
	.B2(\regOut[18][11] ),
	.B1(n572),
	.A2(\regOut[19][11] ),
	.A1(n571), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U1069 (
	.ZN(n832),
	.C2(FE_OFN73_n574),
	.C1(n355),
	.B2(FE_OFN72_n573),
	.B1(n338),
	.A(n835), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U1070 (
	.ZN(n835),
	.B2(\regOut[22][11] ),
	.B1(n577),
	.A2(\regOut[23][11] ),
	.A1(n576), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U1071 (
	.ZN(n831),
	.C2(FE_OFN67_n579),
	.C1(n287),
	.B2(FE_OFN66_n578),
	.B1(n270),
	.A(n836), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U1072 (
	.ZN(n836),
	.B2(\regOut[26][11] ),
	.B1(n582),
	.A2(\regOut[27][11] ),
	.A1(n581), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U1073 (
	.ZN(n830),
	.C2(FE_OFN65_n584),
	.C1(n168),
	.B2(FE_OFN64_n583),
	.B1(n151),
	.A(n837), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U1074 (
	.ZN(n837),
	.B2(\regOut[28][11] ),
	.B1(n587),
	.A2(\regOut[29][11] ),
	.A1(n586), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4_X1 U1075 (
	.ZN(n828),
	.A4(n841),
	.A3(n840),
	.A2(n839),
	.A1(n838), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U1076 (
	.ZN(n841),
	.C2(FE_OFN63_n593),
	.C1(n559),
	.B2(FE_OFN62_n592),
	.B1(n372),
	.A(n842), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U1077 (
	.ZN(n842),
	.B2(\regOut[2][11] ),
	.B1(n596),
	.A2(\regOut[3][11] ),
	.A1(n595), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U1078 (
	.ZN(n840),
	.C2(FE_OFN61_n598),
	.C1(n117),
	.B2(FE_OFN60_n597),
	.B1(n100),
	.A(n843), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U1079 (
	.ZN(n843),
	.B2(\regOut[6][11] ),
	.B1(n601),
	.A2(\regOut[7][11] ),
	.A1(n600), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U1080 (
	.ZN(n839),
	.C2(FE_OFN71_n603),
	.C1(n49),
	.B2(FE_OFN70_n602),
	.B1(n30),
	.A(n844), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U1081 (
	.ZN(n844),
	.B2(\regOut[10][11] ),
	.B1(n606),
	.A2(\regOut[11][11] ),
	.A1(n605), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U1082 (
	.ZN(n838),
	.C2(FE_OFN69_n608),
	.C1(n508),
	.B2(FE_OFN68_n607),
	.B1(n491),
	.A(n845), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U1083 (
	.ZN(n845),
	.B2(\regOut[14][11] ),
	.B1(n611),
	.A2(\regOut[15][11] ),
	.A1(n610), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U1084 (
	.ZN(outB[10]),
	.A2(n847),
	.A1(n846), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4_X1 U1085 (
	.ZN(n847),
	.A4(n851),
	.A3(n850),
	.A2(n849),
	.A1(n848), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U1086 (
	.ZN(n851),
	.C2(FE_OFN75_n569),
	.C1(n441),
	.B2(FE_OFN74_n568),
	.B1(n424),
	.A(n852), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U1087 (
	.ZN(n852),
	.B2(\regOut[18][10] ),
	.B1(n572),
	.A2(\regOut[19][10] ),
	.A1(n571), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U1088 (
	.ZN(n850),
	.C2(FE_OFN73_n574),
	.C1(n356),
	.B2(FE_OFN72_n573),
	.B1(n339),
	.A(n853), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U1089 (
	.ZN(n853),
	.B2(\regOut[22][10] ),
	.B1(n577),
	.A2(\regOut[23][10] ),
	.A1(n576), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U1090 (
	.ZN(n849),
	.C2(FE_OFN67_n579),
	.C1(n288),
	.B2(FE_OFN66_n578),
	.B1(n271),
	.A(n854), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U1091 (
	.ZN(n854),
	.B2(\regOut[26][10] ),
	.B1(n582),
	.A2(\regOut[27][10] ),
	.A1(n581), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U1092 (
	.ZN(n848),
	.C2(FE_OFN65_n584),
	.C1(n169),
	.B2(FE_OFN64_n583),
	.B1(n152),
	.A(n855), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U1093 (
	.ZN(n855),
	.B2(\regOut[28][10] ),
	.B1(n587),
	.A2(\regOut[29][10] ),
	.A1(n586), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4_X1 U1094 (
	.ZN(n846),
	.A4(n859),
	.A3(n858),
	.A2(n857),
	.A1(n856), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U1095 (
	.ZN(n859),
	.C2(FE_OFN63_n593),
	.C1(n560),
	.B2(FE_OFN62_n592),
	.B1(n373),
	.A(n860), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U1096 (
	.ZN(n860),
	.B2(\regOut[2][10] ),
	.B1(n596),
	.A2(\regOut[3][10] ),
	.A1(n595), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U1097 (
	.ZN(n858),
	.C2(FE_OFN61_n598),
	.C1(n118),
	.B2(FE_OFN60_n597),
	.B1(n101),
	.A(n861), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U1098 (
	.ZN(n861),
	.B2(\regOut[6][10] ),
	.B1(n601),
	.A2(\regOut[7][10] ),
	.A1(n600), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U1099 (
	.ZN(n857),
	.C2(FE_OFN71_n603),
	.C1(n50),
	.B2(FE_OFN70_n602),
	.B1(n32),
	.A(n862), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U1100 (
	.ZN(n862),
	.B2(\regOut[10][10] ),
	.B1(n606),
	.A2(\regOut[11][10] ),
	.A1(n605), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U1101 (
	.ZN(n856),
	.C2(FE_OFN69_n608),
	.C1(n509),
	.B2(FE_OFN68_n607),
	.B1(n492),
	.A(n863), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U1102 (
	.ZN(n863),
	.B2(\regOut[14][10] ),
	.B1(n611),
	.A2(\regOut[15][10] ),
	.A1(n610), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U1103 (
	.ZN(outB[0]),
	.A2(n865),
	.A1(n864), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4_X1 U1104 (
	.ZN(n865),
	.A4(n869),
	.A3(n868),
	.A2(n867),
	.A1(n866), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U1105 (
	.ZN(n869),
	.C2(FE_OFN75_n569),
	.C1(n442),
	.B2(FE_OFN74_n568),
	.B1(n425),
	.A(n870), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U1106 (
	.ZN(n870),
	.B2(\regOut[18][0] ),
	.B1(n572),
	.A2(\regOut[19][0] ),
	.A1(n571), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2_X1 U1107 (
	.ZN(n572),
	.A2(n872),
	.A1(n871), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2_X1 U1108 (
	.ZN(n571),
	.A2(n872),
	.A1(n873), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U1109 (
	.ZN(n569),
	.A2(n874),
	.A1(n871), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U1110 (
	.ZN(n568),
	.A2(n874),
	.A1(n873), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U1111 (
	.ZN(n868),
	.C2(FE_OFN73_n574),
	.C1(n357),
	.B2(FE_OFN72_n573),
	.B1(n340),
	.A(n875), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U1112 (
	.ZN(n875),
	.B2(\regOut[22][0] ),
	.B1(n577),
	.A2(\regOut[23][0] ),
	.A1(n576), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2_X1 U1113 (
	.ZN(n577),
	.A2(n876),
	.A1(n871), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2_X1 U1114 (
	.ZN(n576),
	.A2(n876),
	.A1(n873), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U1115 (
	.ZN(n574),
	.A2(n877),
	.A1(n871), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2_X1 U1116 (
	.ZN(n871),
	.A2(n879),
	.A1(n878), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U1117 (
	.ZN(n573),
	.A2(n877),
	.A1(n873), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2_X1 U1118 (
	.ZN(n873),
	.A2(addressB[0]),
	.A1(n878), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2_X1 U1119 (
	.ZN(n878),
	.A2(n880),
	.A1(addressB[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U1120 (
	.ZN(n867),
	.C2(FE_OFN67_n579),
	.C1(n289),
	.B2(FE_OFN66_n578),
	.B1(n272),
	.A(n881), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U1121 (
	.ZN(n881),
	.B2(\regOut[26][0] ),
	.B1(n582),
	.A2(\regOut[27][0] ),
	.A1(n581), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2_X1 U1122 (
	.ZN(n582),
	.A2(n882),
	.A1(n872), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2_X1 U1123 (
	.ZN(n581),
	.A2(n883),
	.A1(n872), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U1124 (
	.ZN(n579),
	.A2(n882),
	.A1(n874), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U1125 (
	.ZN(n578),
	.A2(n883),
	.A1(n874), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U1126 (
	.ZN(n866),
	.C2(FE_OFN65_n584),
	.C1(n170),
	.B2(FE_OFN64_n583),
	.B1(n153),
	.A(n884), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U1127 (
	.ZN(n884),
	.B2(\regOut[28][0] ),
	.B1(n587),
	.A2(\regOut[29][0] ),
	.A1(n586), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2_X1 U1128 (
	.ZN(n587),
	.A2(n882),
	.A1(n877), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2_X1 U1129 (
	.ZN(n586),
	.A2(n883),
	.A1(n877), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U1130 (
	.ZN(n584),
	.A2(n876),
	.A1(n882), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2_X1 U1131 (
	.ZN(n882),
	.A2(n879),
	.A1(n885), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U1132 (
	.ZN(n583),
	.A2(n883),
	.A1(n876), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2_X1 U1133 (
	.ZN(n883),
	.A2(n885),
	.A1(addressB[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2_X1 U1134 (
	.ZN(n885),
	.A2(addressB[3]),
	.A1(addressB[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4_X1 U1135 (
	.ZN(n864),
	.A4(n889),
	.A3(n888),
	.A2(n887),
	.A1(n886), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U1136 (
	.ZN(n889),
	.C2(FE_OFN63_n593),
	.C1(n561),
	.B2(FE_OFN62_n592),
	.B1(n374),
	.A(n890), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U1137 (
	.ZN(n890),
	.B2(\regOut[2][0] ),
	.B1(n596),
	.A2(\regOut[3][0] ),
	.A1(n595), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2_X1 U1138 (
	.ZN(n596),
	.A2(n872),
	.A1(n891), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2_X1 U1139 (
	.ZN(n595),
	.A2(n872),
	.A1(n892), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U1140 (
	.ZN(n593),
	.A2(n874),
	.A1(n891), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U1141 (
	.ZN(n592),
	.A2(n874),
	.A1(n892), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U1142 (
	.ZN(n888),
	.C2(FE_OFN61_n598),
	.C1(n119),
	.B2(FE_OFN60_n597),
	.B1(n102),
	.A(n893), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U1143 (
	.ZN(n893),
	.B2(\regOut[6][0] ),
	.B1(n601),
	.A2(\regOut[7][0] ),
	.A1(n600), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2_X1 U1144 (
	.ZN(n601),
	.A2(n876),
	.A1(n891), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2_X1 U1145 (
	.ZN(n600),
	.A2(n876),
	.A1(n892), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U1146 (
	.ZN(n598),
	.A2(n877),
	.A1(n891), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2_X1 U1147 (
	.ZN(n891),
	.A2(n879),
	.A1(n894), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U1148 (
	.ZN(n597),
	.A2(n877),
	.A1(n892), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2_X1 U1149 (
	.ZN(n892),
	.A2(addressB[0]),
	.A1(n894), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2_X1 U1150 (
	.ZN(n894),
	.A2(addressB[4]),
	.A1(addressB[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U1151 (
	.ZN(n887),
	.C2(FE_OFN71_n603),
	.C1(n51),
	.B2(FE_OFN70_n602),
	.B1(n34),
	.A(n895), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U1152 (
	.ZN(n895),
	.B2(\regOut[10][0] ),
	.B1(n606),
	.A2(\regOut[11][0] ),
	.A1(n605), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2_X1 U1153 (
	.ZN(n606),
	.A2(n872),
	.A1(n896), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2_X1 U1154 (
	.ZN(n605),
	.A2(n872),
	.A1(n897), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2_X1 U1155 (
	.ZN(n872),
	.A2(addressB[2]),
	.A1(n898), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U1156 (
	.ZN(n603),
	.A2(n874),
	.A1(n896), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U1157 (
	.ZN(n602),
	.A2(n874),
	.A1(n897), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2_X2 U1158 (
	.ZN(n874),
	.A2(addressB[2]),
	.A1(addressB[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U1159 (
	.ZN(n886),
	.C2(FE_OFN69_n608),
	.C1(n510),
	.B2(FE_OFN68_n607),
	.B1(n493),
	.A(n899), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U1160 (
	.ZN(n899),
	.B2(\regOut[14][0] ),
	.B1(n611),
	.A2(\regOut[15][0] ),
	.A1(n610), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2_X1 U1161 (
	.ZN(n611),
	.A2(n876),
	.A1(n896), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2_X1 U1162 (
	.ZN(n610),
	.A2(n876),
	.A1(n897), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2_X1 U1163 (
	.ZN(n876),
	.A2(n898),
	.A1(n900), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1164 (
	.ZN(n898),
	.A(addressB[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U1165 (
	.ZN(n608),
	.A2(n877),
	.A1(n896), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2_X1 U1166 (
	.ZN(n896),
	.A2(n879),
	.A1(n901), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1167 (
	.ZN(n879),
	.A(addressB[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U1168 (
	.ZN(n607),
	.A2(n877),
	.A1(n897), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2_X2 U1169 (
	.ZN(n877),
	.A2(addressB[1]),
	.A1(n900), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1170 (
	.ZN(n900),
	.A(addressB[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2_X1 U1171 (
	.ZN(n897),
	.A2(addressB[0]),
	.A1(n901), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2_X1 U1172 (
	.ZN(n901),
	.A2(addressB[4]),
	.A1(n880), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1173 (
	.ZN(n880),
	.A(addressB[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U1174 (
	.ZN(outA[9]),
	.A2(n903),
	.A1(n902), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4_X1 U1175 (
	.ZN(n903),
	.A4(n907),
	.A3(n906),
	.A2(n905),
	.A1(n904), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U1176 (
	.ZN(n907),
	.C2(n909),
	.C1(n427),
	.B2(n908),
	.B1(n410),
	.A(n910), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U1177 (
	.ZN(n910),
	.B2(\regOut[18][9] ),
	.B1(n912),
	.A2(\regOut[19][9] ),
	.A1(n911), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1178 (
	.ZN(n427),
	.A(\regOut[16][9] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1179 (
	.ZN(n410),
	.A(\regOut[17][9] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U1180 (
	.ZN(n906),
	.C2(n914),
	.C1(n342),
	.B2(n913),
	.B1(n325),
	.A(n915), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U1181 (
	.ZN(n915),
	.B2(\regOut[22][9] ),
	.B1(n917),
	.A2(\regOut[23][9] ),
	.A1(n916), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1182 (
	.ZN(n342),
	.A(\regOut[20][9] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1183 (
	.ZN(n325),
	.A(\regOut[21][9] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U1184 (
	.ZN(n905),
	.C2(n919),
	.C1(n274),
	.B2(n918),
	.B1(n257),
	.A(n920), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U1185 (
	.ZN(n920),
	.B2(\regOut[26][9] ),
	.B1(n922),
	.A2(\regOut[27][9] ),
	.A1(n921), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1186 (
	.ZN(n274),
	.A(\regOut[24][9] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1187 (
	.ZN(n257),
	.A(\regOut[25][9] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U1188 (
	.ZN(n904),
	.C2(n924),
	.C1(n155),
	.B2(n923),
	.B1(n138),
	.A(n925), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U1189 (
	.ZN(n925),
	.B2(\regOut[28][9] ),
	.B1(n927),
	.A2(\regOut[29][9] ),
	.A1(n926), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1190 (
	.ZN(n155),
	.A(\regOut[30][9] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1191 (
	.ZN(n138),
	.A(\regOut[31][9] ), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4_X1 U1192 (
	.ZN(n902),
	.A4(n931),
	.A3(n930),
	.A2(n929),
	.A1(n928), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U1193 (
	.ZN(n931),
	.C2(n933),
	.C1(n546),
	.B2(n932),
	.B1(n359),
	.A(n934), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U1194 (
	.ZN(n934),
	.B2(\regOut[2][9] ),
	.B1(n936),
	.A2(\regOut[3][9] ),
	.A1(n935), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1195 (
	.ZN(n546),
	.A(\regOut[0][9] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1196 (
	.ZN(n359),
	.A(\regOut[1][9] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U1197 (
	.ZN(n930),
	.C2(n938),
	.C1(n104),
	.B2(n937),
	.B1(n87),
	.A(n939), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U1198 (
	.ZN(n939),
	.B2(\regOut[6][9] ),
	.B1(n941),
	.A2(\regOut[7][9] ),
	.A1(n940), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1199 (
	.ZN(n104),
	.A(\regOut[4][9] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1200 (
	.ZN(n87),
	.A(\regOut[5][9] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U1201 (
	.ZN(n929),
	.C2(n943),
	.C1(n36),
	.B2(n942),
	.B1(n4),
	.A(n944), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U1202 (
	.ZN(n944),
	.B2(\regOut[10][9] ),
	.B1(n946),
	.A2(\regOut[11][9] ),
	.A1(n945), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1203 (
	.ZN(n36),
	.A(\regOut[8][9] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1204 (
	.ZN(n4),
	.A(\regOut[9][9] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U1205 (
	.ZN(n928),
	.C2(n948),
	.C1(n495),
	.B2(n947),
	.B1(n478),
	.A(n949), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U1206 (
	.ZN(n949),
	.B2(\regOut[14][9] ),
	.B1(n951),
	.A2(\regOut[15][9] ),
	.A1(n950), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1207 (
	.ZN(n495),
	.A(\regOut[12][9] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1208 (
	.ZN(n478),
	.A(\regOut[13][9] ), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U1209 (
	.ZN(outA[8]),
	.A2(n953),
	.A1(n952), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4_X1 U1210 (
	.ZN(n953),
	.A4(n957),
	.A3(n956),
	.A2(n955),
	.A1(n954), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U1211 (
	.ZN(n957),
	.C2(n909),
	.C1(n428),
	.B2(n908),
	.B1(n411),
	.A(n958), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U1212 (
	.ZN(n958),
	.B2(\regOut[18][8] ),
	.B1(n912),
	.A2(\regOut[19][8] ),
	.A1(n911), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1213 (
	.ZN(n428),
	.A(\regOut[16][8] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1214 (
	.ZN(n411),
	.A(\regOut[17][8] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U1215 (
	.ZN(n956),
	.C2(n914),
	.C1(n343),
	.B2(n913),
	.B1(n326),
	.A(n959), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U1216 (
	.ZN(n959),
	.B2(\regOut[22][8] ),
	.B1(n917),
	.A2(\regOut[23][8] ),
	.A1(n916), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1217 (
	.ZN(n343),
	.A(\regOut[20][8] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1218 (
	.ZN(n326),
	.A(\regOut[21][8] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U1219 (
	.ZN(n955),
	.C2(n919),
	.C1(n275),
	.B2(n918),
	.B1(n258),
	.A(n960), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U1220 (
	.ZN(n960),
	.B2(\regOut[26][8] ),
	.B1(n922),
	.A2(\regOut[27][8] ),
	.A1(n921), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1221 (
	.ZN(n275),
	.A(\regOut[24][8] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1222 (
	.ZN(n258),
	.A(\regOut[25][8] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U1223 (
	.ZN(n954),
	.C2(n924),
	.C1(n156),
	.B2(n923),
	.B1(n139),
	.A(n961), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U1224 (
	.ZN(n961),
	.B2(\regOut[28][8] ),
	.B1(n927),
	.A2(\regOut[29][8] ),
	.A1(n926), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1225 (
	.ZN(n156),
	.A(\regOut[30][8] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1226 (
	.ZN(n139),
	.A(\regOut[31][8] ), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4_X1 U1227 (
	.ZN(n952),
	.A4(n965),
	.A3(n964),
	.A2(n963),
	.A1(n962), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U1228 (
	.ZN(n965),
	.C2(n933),
	.C1(n547),
	.B2(n932),
	.B1(n360),
	.A(n966), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U1229 (
	.ZN(n966),
	.B2(\regOut[2][8] ),
	.B1(n936),
	.A2(\regOut[3][8] ),
	.A1(n935), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1230 (
	.ZN(n547),
	.A(\regOut[0][8] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1231 (
	.ZN(n360),
	.A(\regOut[1][8] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U1232 (
	.ZN(n964),
	.C2(n938),
	.C1(n105),
	.B2(n937),
	.B1(n88),
	.A(n967), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U1233 (
	.ZN(n967),
	.B2(\regOut[6][8] ),
	.B1(n941),
	.A2(\regOut[7][8] ),
	.A1(n940), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1234 (
	.ZN(n105),
	.A(\regOut[4][8] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1235 (
	.ZN(n88),
	.A(\regOut[5][8] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U1236 (
	.ZN(n963),
	.C2(n943),
	.C1(n37),
	.B2(n942),
	.B1(n6),
	.A(n968), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U1237 (
	.ZN(n968),
	.B2(\regOut[10][8] ),
	.B1(n946),
	.A2(\regOut[11][8] ),
	.A1(n945), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1238 (
	.ZN(n37),
	.A(\regOut[8][8] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1239 (
	.ZN(n6),
	.A(\regOut[9][8] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U1240 (
	.ZN(n962),
	.C2(n948),
	.C1(n496),
	.B2(n947),
	.B1(n479),
	.A(n969), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U1241 (
	.ZN(n969),
	.B2(\regOut[14][8] ),
	.B1(n951),
	.A2(\regOut[15][8] ),
	.A1(n950), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1242 (
	.ZN(n496),
	.A(\regOut[12][8] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1243 (
	.ZN(n479),
	.A(\regOut[13][8] ), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U1244 (
	.ZN(outA[7]),
	.A2(n971),
	.A1(n970), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4_X1 U1245 (
	.ZN(n971),
	.A4(n975),
	.A3(n974),
	.A2(n973),
	.A1(n972), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U1246 (
	.ZN(n975),
	.C2(n909),
	.C1(n429),
	.B2(n908),
	.B1(n412),
	.A(n976), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U1247 (
	.ZN(n976),
	.B2(\regOut[18][7] ),
	.B1(n912),
	.A2(\regOut[19][7] ),
	.A1(n911), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1248 (
	.ZN(n429),
	.A(\regOut[16][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1249 (
	.ZN(n412),
	.A(\regOut[17][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U1250 (
	.ZN(n974),
	.C2(n914),
	.C1(n344),
	.B2(n913),
	.B1(n327),
	.A(n977), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U1251 (
	.ZN(n977),
	.B2(\regOut[22][7] ),
	.B1(n917),
	.A2(\regOut[23][7] ),
	.A1(n916), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1252 (
	.ZN(n344),
	.A(\regOut[20][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1253 (
	.ZN(n327),
	.A(\regOut[21][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U1254 (
	.ZN(n973),
	.C2(n919),
	.C1(n276),
	.B2(n918),
	.B1(n259),
	.A(n978), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U1255 (
	.ZN(n978),
	.B2(\regOut[26][7] ),
	.B1(n922),
	.A2(\regOut[27][7] ),
	.A1(n921), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1256 (
	.ZN(n276),
	.A(\regOut[24][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1257 (
	.ZN(n259),
	.A(\regOut[25][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U1258 (
	.ZN(n972),
	.C2(n924),
	.C1(n157),
	.B2(n923),
	.B1(n140),
	.A(n979), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U1259 (
	.ZN(n979),
	.B2(\regOut[28][7] ),
	.B1(n927),
	.A2(\regOut[29][7] ),
	.A1(n926), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1260 (
	.ZN(n157),
	.A(\regOut[30][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1261 (
	.ZN(n140),
	.A(\regOut[31][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4_X1 U1262 (
	.ZN(n970),
	.A4(n983),
	.A3(n982),
	.A2(n981),
	.A1(n980), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U1263 (
	.ZN(n983),
	.C2(n933),
	.C1(n548),
	.B2(n932),
	.B1(n361),
	.A(n984), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U1264 (
	.ZN(n984),
	.B2(\regOut[2][7] ),
	.B1(n936),
	.A2(\regOut[3][7] ),
	.A1(n935), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1265 (
	.ZN(n548),
	.A(\regOut[0][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1266 (
	.ZN(n361),
	.A(\regOut[1][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U1267 (
	.ZN(n982),
	.C2(n938),
	.C1(n106),
	.B2(n937),
	.B1(n89),
	.A(n985), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U1268 (
	.ZN(n985),
	.B2(\regOut[6][7] ),
	.B1(n941),
	.A2(\regOut[7][7] ),
	.A1(n940), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1269 (
	.ZN(n106),
	.A(\regOut[4][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1270 (
	.ZN(n89),
	.A(\regOut[5][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U1271 (
	.ZN(n981),
	.C2(n943),
	.C1(n38),
	.B2(n942),
	.B1(n8),
	.A(n986), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U1272 (
	.ZN(n986),
	.B2(\regOut[10][7] ),
	.B1(n946),
	.A2(\regOut[11][7] ),
	.A1(n945), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1273 (
	.ZN(n38),
	.A(\regOut[8][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1274 (
	.ZN(n8),
	.A(\regOut[9][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U1275 (
	.ZN(n980),
	.C2(n948),
	.C1(n497),
	.B2(n947),
	.B1(n480),
	.A(n987), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U1276 (
	.ZN(n987),
	.B2(\regOut[14][7] ),
	.B1(n951),
	.A2(\regOut[15][7] ),
	.A1(n950), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1277 (
	.ZN(n497),
	.A(\regOut[12][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1278 (
	.ZN(n480),
	.A(\regOut[13][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U1279 (
	.ZN(outA[6]),
	.A2(n989),
	.A1(n988), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4_X1 U1280 (
	.ZN(n989),
	.A4(n993),
	.A3(n992),
	.A2(n991),
	.A1(n990), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U1281 (
	.ZN(n993),
	.C2(n909),
	.C1(n430),
	.B2(n908),
	.B1(n413),
	.A(n994), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U1282 (
	.ZN(n994),
	.B2(\regOut[18][6] ),
	.B1(n912),
	.A2(\regOut[19][6] ),
	.A1(n911), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1283 (
	.ZN(n430),
	.A(\regOut[16][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1284 (
	.ZN(n413),
	.A(\regOut[17][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U1285 (
	.ZN(n992),
	.C2(n914),
	.C1(n345),
	.B2(n913),
	.B1(n328),
	.A(n995), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U1286 (
	.ZN(n995),
	.B2(\regOut[22][6] ),
	.B1(n917),
	.A2(\regOut[23][6] ),
	.A1(n916), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1287 (
	.ZN(n345),
	.A(\regOut[20][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1288 (
	.ZN(n328),
	.A(\regOut[21][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U1289 (
	.ZN(n991),
	.C2(n919),
	.C1(n277),
	.B2(n918),
	.B1(n260),
	.A(n996), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U1290 (
	.ZN(n996),
	.B2(\regOut[26][6] ),
	.B1(n922),
	.A2(\regOut[27][6] ),
	.A1(n921), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1291 (
	.ZN(n277),
	.A(\regOut[24][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1292 (
	.ZN(n260),
	.A(\regOut[25][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U1293 (
	.ZN(n990),
	.C2(n924),
	.C1(n158),
	.B2(n923),
	.B1(n141),
	.A(n997), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U1294 (
	.ZN(n997),
	.B2(\regOut[28][6] ),
	.B1(n927),
	.A2(\regOut[29][6] ),
	.A1(n926), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1295 (
	.ZN(n158),
	.A(\regOut[30][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1296 (
	.ZN(n141),
	.A(\regOut[31][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4_X1 U1297 (
	.ZN(n988),
	.A4(n1001),
	.A3(n1000),
	.A2(n999),
	.A1(n998), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U1298 (
	.ZN(n1001),
	.C2(n933),
	.C1(n549),
	.B2(n932),
	.B1(n362),
	.A(n1002), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U1299 (
	.ZN(n1002),
	.B2(\regOut[2][6] ),
	.B1(n936),
	.A2(\regOut[3][6] ),
	.A1(n935), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1300 (
	.ZN(n549),
	.A(\regOut[0][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1301 (
	.ZN(n362),
	.A(\regOut[1][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U1302 (
	.ZN(n1000),
	.C2(n938),
	.C1(n107),
	.B2(n937),
	.B1(n90),
	.A(n1003), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U1303 (
	.ZN(n1003),
	.B2(\regOut[6][6] ),
	.B1(n941),
	.A2(\regOut[7][6] ),
	.A1(n940), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1304 (
	.ZN(n107),
	.A(\regOut[4][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1305 (
	.ZN(n90),
	.A(\regOut[5][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U1306 (
	.ZN(n999),
	.C2(n943),
	.C1(n39),
	.B2(n942),
	.B1(n10),
	.A(n1004), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U1307 (
	.ZN(n1004),
	.B2(\regOut[10][6] ),
	.B1(n946),
	.A2(\regOut[11][6] ),
	.A1(n945), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1308 (
	.ZN(n39),
	.A(\regOut[8][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1309 (
	.ZN(n10),
	.A(\regOut[9][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U1310 (
	.ZN(n998),
	.C2(n948),
	.C1(n498),
	.B2(n947),
	.B1(n481),
	.A(n1005), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U1311 (
	.ZN(n1005),
	.B2(\regOut[14][6] ),
	.B1(n951),
	.A2(\regOut[15][6] ),
	.A1(n950), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1312 (
	.ZN(n498),
	.A(\regOut[12][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1313 (
	.ZN(n481),
	.A(\regOut[13][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U1314 (
	.ZN(outA[5]),
	.A2(n1007),
	.A1(n1006), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4_X1 U1315 (
	.ZN(n1007),
	.A4(n1011),
	.A3(n1010),
	.A2(n1009),
	.A1(n1008), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U1316 (
	.ZN(n1011),
	.C2(n909),
	.C1(n431),
	.B2(n908),
	.B1(n414),
	.A(n1012), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U1317 (
	.ZN(n1012),
	.B2(\regOut[18][5] ),
	.B1(n912),
	.A2(\regOut[19][5] ),
	.A1(n911), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1318 (
	.ZN(n431),
	.A(\regOut[16][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1319 (
	.ZN(n414),
	.A(\regOut[17][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U1320 (
	.ZN(n1010),
	.C2(n914),
	.C1(n346),
	.B2(n913),
	.B1(n329),
	.A(n1013), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U1321 (
	.ZN(n1013),
	.B2(\regOut[22][5] ),
	.B1(n917),
	.A2(\regOut[23][5] ),
	.A1(n916), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1322 (
	.ZN(n346),
	.A(\regOut[20][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1323 (
	.ZN(n329),
	.A(\regOut[21][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U1324 (
	.ZN(n1009),
	.C2(n919),
	.C1(n278),
	.B2(n918),
	.B1(n261),
	.A(n1014), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U1325 (
	.ZN(n1014),
	.B2(\regOut[26][5] ),
	.B1(n922),
	.A2(\regOut[27][5] ),
	.A1(n921), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1326 (
	.ZN(n278),
	.A(\regOut[24][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1327 (
	.ZN(n261),
	.A(\regOut[25][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U1328 (
	.ZN(n1008),
	.C2(n924),
	.C1(n159),
	.B2(n923),
	.B1(n142),
	.A(n1015), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U1329 (
	.ZN(n1015),
	.B2(\regOut[28][5] ),
	.B1(n927),
	.A2(\regOut[29][5] ),
	.A1(n926), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1330 (
	.ZN(n159),
	.A(\regOut[30][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1331 (
	.ZN(n142),
	.A(\regOut[31][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4_X1 U1332 (
	.ZN(n1006),
	.A4(n1019),
	.A3(n1018),
	.A2(n1017),
	.A1(n1016), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U1333 (
	.ZN(n1019),
	.C2(n933),
	.C1(n550),
	.B2(n932),
	.B1(n363),
	.A(n1020), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U1334 (
	.ZN(n1020),
	.B2(\regOut[2][5] ),
	.B1(n936),
	.A2(\regOut[3][5] ),
	.A1(n935), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1335 (
	.ZN(n550),
	.A(\regOut[0][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1336 (
	.ZN(n363),
	.A(\regOut[1][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U1337 (
	.ZN(n1018),
	.C2(n938),
	.C1(n108),
	.B2(n937),
	.B1(n91),
	.A(n1021), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U1338 (
	.ZN(n1021),
	.B2(\regOut[6][5] ),
	.B1(n941),
	.A2(\regOut[7][5] ),
	.A1(n940), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1339 (
	.ZN(n108),
	.A(\regOut[4][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1340 (
	.ZN(n91),
	.A(\regOut[5][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U1341 (
	.ZN(n1017),
	.C2(n943),
	.C1(n40),
	.B2(n942),
	.B1(n12),
	.A(n1022), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U1342 (
	.ZN(n1022),
	.B2(\regOut[10][5] ),
	.B1(n946),
	.A2(\regOut[11][5] ),
	.A1(n945), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1343 (
	.ZN(n40),
	.A(\regOut[8][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1344 (
	.ZN(n12),
	.A(\regOut[9][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U1345 (
	.ZN(n1016),
	.C2(n948),
	.C1(n499),
	.B2(n947),
	.B1(n482),
	.A(n1023), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U1346 (
	.ZN(n1023),
	.B2(\regOut[14][5] ),
	.B1(n951),
	.A2(\regOut[15][5] ),
	.A1(n950), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1347 (
	.ZN(n499),
	.A(\regOut[12][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1348 (
	.ZN(n482),
	.A(\regOut[13][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U1349 (
	.ZN(outA[4]),
	.A2(n1025),
	.A1(n1024), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4_X1 U1350 (
	.ZN(n1025),
	.A4(n1029),
	.A3(n1028),
	.A2(n1027),
	.A1(n1026), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U1351 (
	.ZN(n1029),
	.C2(n909),
	.C1(n432),
	.B2(n908),
	.B1(n415),
	.A(n1030), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U1352 (
	.ZN(n1030),
	.B2(\regOut[18][4] ),
	.B1(n912),
	.A2(\regOut[19][4] ),
	.A1(n911), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1353 (
	.ZN(n432),
	.A(\regOut[16][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1354 (
	.ZN(n415),
	.A(\regOut[17][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U1355 (
	.ZN(n1028),
	.C2(n914),
	.C1(n347),
	.B2(n913),
	.B1(n330),
	.A(n1031), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U1356 (
	.ZN(n1031),
	.B2(\regOut[22][4] ),
	.B1(n917),
	.A2(\regOut[23][4] ),
	.A1(n916), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1357 (
	.ZN(n347),
	.A(\regOut[20][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1358 (
	.ZN(n330),
	.A(\regOut[21][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U1359 (
	.ZN(n1027),
	.C2(n919),
	.C1(n279),
	.B2(n918),
	.B1(n262),
	.A(n1032), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U1360 (
	.ZN(n1032),
	.B2(\regOut[26][4] ),
	.B1(n922),
	.A2(\regOut[27][4] ),
	.A1(n921), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1361 (
	.ZN(n279),
	.A(\regOut[24][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1362 (
	.ZN(n262),
	.A(\regOut[25][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U1363 (
	.ZN(n1026),
	.C2(n924),
	.C1(n160),
	.B2(n923),
	.B1(n143),
	.A(n1033), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U1364 (
	.ZN(n1033),
	.B2(\regOut[28][4] ),
	.B1(n927),
	.A2(\regOut[29][4] ),
	.A1(n926), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1365 (
	.ZN(n160),
	.A(\regOut[30][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1366 (
	.ZN(n143),
	.A(\regOut[31][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4_X1 U1367 (
	.ZN(n1024),
	.A4(n1037),
	.A3(n1036),
	.A2(n1035),
	.A1(n1034), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U1368 (
	.ZN(n1037),
	.C2(n933),
	.C1(n551),
	.B2(n932),
	.B1(n364),
	.A(n1038), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U1369 (
	.ZN(n1038),
	.B2(\regOut[2][4] ),
	.B1(n936),
	.A2(\regOut[3][4] ),
	.A1(n935), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1370 (
	.ZN(n551),
	.A(\regOut[0][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1371 (
	.ZN(n364),
	.A(\regOut[1][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U1372 (
	.ZN(n1036),
	.C2(n938),
	.C1(n109),
	.B2(n937),
	.B1(n92),
	.A(n1039), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U1373 (
	.ZN(n1039),
	.B2(\regOut[6][4] ),
	.B1(n941),
	.A2(\regOut[7][4] ),
	.A1(n940), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1374 (
	.ZN(n109),
	.A(\regOut[4][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1375 (
	.ZN(n92),
	.A(\regOut[5][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U1376 (
	.ZN(n1035),
	.C2(n943),
	.C1(n41),
	.B2(n942),
	.B1(n14),
	.A(n1040), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U1377 (
	.ZN(n1040),
	.B2(\regOut[10][4] ),
	.B1(n946),
	.A2(\regOut[11][4] ),
	.A1(n945), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1378 (
	.ZN(n41),
	.A(\regOut[8][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1379 (
	.ZN(n14),
	.A(\regOut[9][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U1380 (
	.ZN(n1034),
	.C2(n948),
	.C1(n500),
	.B2(n947),
	.B1(n483),
	.A(n1041), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U1381 (
	.ZN(n1041),
	.B2(\regOut[14][4] ),
	.B1(n951),
	.A2(\regOut[15][4] ),
	.A1(n950), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1382 (
	.ZN(n500),
	.A(\regOut[12][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1383 (
	.ZN(n483),
	.A(\regOut[13][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U1384 (
	.ZN(outA[3]),
	.A2(n1043),
	.A1(n1042), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4_X1 U1385 (
	.ZN(n1043),
	.A4(n1047),
	.A3(n1046),
	.A2(n1045),
	.A1(n1044), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U1386 (
	.ZN(n1047),
	.C2(n909),
	.C1(n433),
	.B2(n908),
	.B1(n416),
	.A(n1048), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U1387 (
	.ZN(n1048),
	.B2(\regOut[18][3] ),
	.B1(n912),
	.A2(\regOut[19][3] ),
	.A1(n911), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1388 (
	.ZN(n433),
	.A(\regOut[16][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1389 (
	.ZN(n416),
	.A(\regOut[17][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U1390 (
	.ZN(n1046),
	.C2(n914),
	.C1(n348),
	.B2(n913),
	.B1(n331),
	.A(n1049), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U1391 (
	.ZN(n1049),
	.B2(\regOut[22][3] ),
	.B1(n917),
	.A2(\regOut[23][3] ),
	.A1(n916), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1392 (
	.ZN(n348),
	.A(\regOut[20][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1393 (
	.ZN(n331),
	.A(\regOut[21][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U1394 (
	.ZN(n1045),
	.C2(n919),
	.C1(n280),
	.B2(n918),
	.B1(n263),
	.A(n1050), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U1395 (
	.ZN(n1050),
	.B2(\regOut[26][3] ),
	.B1(n922),
	.A2(\regOut[27][3] ),
	.A1(n921), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1396 (
	.ZN(n280),
	.A(\regOut[24][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1397 (
	.ZN(n263),
	.A(\regOut[25][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U1398 (
	.ZN(n1044),
	.C2(n924),
	.C1(n161),
	.B2(n923),
	.B1(n144),
	.A(n1051), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U1399 (
	.ZN(n1051),
	.B2(\regOut[28][3] ),
	.B1(n927),
	.A2(\regOut[29][3] ),
	.A1(n926), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1400 (
	.ZN(n161),
	.A(\regOut[30][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1401 (
	.ZN(n144),
	.A(\regOut[31][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4_X1 U1402 (
	.ZN(n1042),
	.A4(n1055),
	.A3(n1054),
	.A2(n1053),
	.A1(n1052), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U1403 (
	.ZN(n1055),
	.C2(n933),
	.C1(n552),
	.B2(n932),
	.B1(n365),
	.A(n1056), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U1404 (
	.ZN(n1056),
	.B2(\regOut[2][3] ),
	.B1(n936),
	.A2(\regOut[3][3] ),
	.A1(n935), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1405 (
	.ZN(n552),
	.A(\regOut[0][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1406 (
	.ZN(n365),
	.A(\regOut[1][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U1407 (
	.ZN(n1054),
	.C2(n938),
	.C1(n110),
	.B2(n937),
	.B1(n93),
	.A(n1057), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U1408 (
	.ZN(n1057),
	.B2(\regOut[6][3] ),
	.B1(n941),
	.A2(\regOut[7][3] ),
	.A1(n940), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1409 (
	.ZN(n110),
	.A(\regOut[4][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1410 (
	.ZN(n93),
	.A(\regOut[5][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U1411 (
	.ZN(n1053),
	.C2(n943),
	.C1(n42),
	.B2(n942),
	.B1(n16),
	.A(n1058), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U1412 (
	.ZN(n1058),
	.B2(\regOut[10][3] ),
	.B1(n946),
	.A2(\regOut[11][3] ),
	.A1(n945), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1413 (
	.ZN(n42),
	.A(\regOut[8][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1414 (
	.ZN(n16),
	.A(\regOut[9][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U1415 (
	.ZN(n1052),
	.C2(n948),
	.C1(n501),
	.B2(n947),
	.B1(n484),
	.A(n1059), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U1416 (
	.ZN(n1059),
	.B2(\regOut[14][3] ),
	.B1(n951),
	.A2(\regOut[15][3] ),
	.A1(n950), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1417 (
	.ZN(n501),
	.A(\regOut[12][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1418 (
	.ZN(n484),
	.A(\regOut[13][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U1419 (
	.ZN(outA[2]),
	.A2(n1061),
	.A1(n1060), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4_X1 U1420 (
	.ZN(n1061),
	.A4(n1065),
	.A3(n1064),
	.A2(n1063),
	.A1(n1062), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U1421 (
	.ZN(n1065),
	.C2(n909),
	.C1(n434),
	.B2(n908),
	.B1(n417),
	.A(n1066), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U1422 (
	.ZN(n1066),
	.B2(\regOut[18][2] ),
	.B1(n912),
	.A2(\regOut[19][2] ),
	.A1(n911), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1423 (
	.ZN(n434),
	.A(\regOut[16][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1424 (
	.ZN(n417),
	.A(\regOut[17][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U1425 (
	.ZN(n1064),
	.C2(n914),
	.C1(n349),
	.B2(n913),
	.B1(n332),
	.A(n1067), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U1426 (
	.ZN(n1067),
	.B2(\regOut[22][2] ),
	.B1(n917),
	.A2(\regOut[23][2] ),
	.A1(n916), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1427 (
	.ZN(n349),
	.A(\regOut[20][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1428 (
	.ZN(n332),
	.A(\regOut[21][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U1429 (
	.ZN(n1063),
	.C2(n919),
	.C1(n281),
	.B2(n918),
	.B1(n264),
	.A(n1068), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U1430 (
	.ZN(n1068),
	.B2(\regOut[26][2] ),
	.B1(n922),
	.A2(\regOut[27][2] ),
	.A1(n921), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1431 (
	.ZN(n281),
	.A(\regOut[24][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1432 (
	.ZN(n264),
	.A(\regOut[25][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U1433 (
	.ZN(n1062),
	.C2(n924),
	.C1(n162),
	.B2(n923),
	.B1(n145),
	.A(n1069), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U1434 (
	.ZN(n1069),
	.B2(\regOut[28][2] ),
	.B1(n927),
	.A2(\regOut[29][2] ),
	.A1(n926), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1435 (
	.ZN(n162),
	.A(\regOut[30][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1436 (
	.ZN(n145),
	.A(\regOut[31][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4_X1 U1437 (
	.ZN(n1060),
	.A4(n1073),
	.A3(n1072),
	.A2(n1071),
	.A1(n1070), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U1438 (
	.ZN(n1073),
	.C2(n933),
	.C1(n553),
	.B2(n932),
	.B1(n366),
	.A(n1074), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U1439 (
	.ZN(n1074),
	.B2(\regOut[2][2] ),
	.B1(n936),
	.A2(\regOut[3][2] ),
	.A1(n935), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1440 (
	.ZN(n553),
	.A(\regOut[0][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1441 (
	.ZN(n366),
	.A(\regOut[1][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U1442 (
	.ZN(n1072),
	.C2(n938),
	.C1(n111),
	.B2(n937),
	.B1(n94),
	.A(n1075), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U1443 (
	.ZN(n1075),
	.B2(\regOut[6][2] ),
	.B1(n941),
	.A2(\regOut[7][2] ),
	.A1(n940), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1444 (
	.ZN(n111),
	.A(\regOut[4][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1445 (
	.ZN(n94),
	.A(\regOut[5][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U1446 (
	.ZN(n1071),
	.C2(n943),
	.C1(n43),
	.B2(n942),
	.B1(n18),
	.A(n1076), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U1447 (
	.ZN(n1076),
	.B2(\regOut[10][2] ),
	.B1(n946),
	.A2(\regOut[11][2] ),
	.A1(n945), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1448 (
	.ZN(n43),
	.A(\regOut[8][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1449 (
	.ZN(n18),
	.A(\regOut[9][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U1450 (
	.ZN(n1070),
	.C2(n948),
	.C1(n502),
	.B2(n947),
	.B1(n485),
	.A(n1077), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U1451 (
	.ZN(n1077),
	.B2(\regOut[14][2] ),
	.B1(n951),
	.A2(\regOut[15][2] ),
	.A1(n950), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1452 (
	.ZN(n502),
	.A(\regOut[12][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1453 (
	.ZN(n485),
	.A(\regOut[13][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U1454 (
	.ZN(outA[1]),
	.A2(n1079),
	.A1(n1078), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4_X1 U1455 (
	.ZN(n1079),
	.A4(n1083),
	.A3(n1082),
	.A2(n1081),
	.A1(n1080), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U1456 (
	.ZN(n1083),
	.C2(n909),
	.C1(n435),
	.B2(n908),
	.B1(n418),
	.A(n1084), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U1457 (
	.ZN(n1084),
	.B2(\regOut[18][1] ),
	.B1(n912),
	.A2(\regOut[19][1] ),
	.A1(n911), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1458 (
	.ZN(n435),
	.A(\regOut[16][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1459 (
	.ZN(n418),
	.A(\regOut[17][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U1460 (
	.ZN(n1082),
	.C2(n914),
	.C1(n350),
	.B2(n913),
	.B1(n333),
	.A(n1085), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U1461 (
	.ZN(n1085),
	.B2(\regOut[22][1] ),
	.B1(n917),
	.A2(\regOut[23][1] ),
	.A1(n916), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1462 (
	.ZN(n350),
	.A(\regOut[20][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1463 (
	.ZN(n333),
	.A(\regOut[21][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U1464 (
	.ZN(n1081),
	.C2(n919),
	.C1(n282),
	.B2(n918),
	.B1(n265),
	.A(n1086), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U1465 (
	.ZN(n1086),
	.B2(\regOut[26][1] ),
	.B1(n922),
	.A2(\regOut[27][1] ),
	.A1(n921), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1466 (
	.ZN(n282),
	.A(\regOut[24][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1467 (
	.ZN(n265),
	.A(\regOut[25][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U1468 (
	.ZN(n1080),
	.C2(n924),
	.C1(n163),
	.B2(n923),
	.B1(n146),
	.A(n1087), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U1469 (
	.ZN(n1087),
	.B2(\regOut[28][1] ),
	.B1(n927),
	.A2(\regOut[29][1] ),
	.A1(n926), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1470 (
	.ZN(n163),
	.A(\regOut[30][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1471 (
	.ZN(n146),
	.A(\regOut[31][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4_X1 U1472 (
	.ZN(n1078),
	.A4(n1091),
	.A3(n1090),
	.A2(n1089),
	.A1(n1088), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U1473 (
	.ZN(n1091),
	.C2(n933),
	.C1(n554),
	.B2(n932),
	.B1(n367),
	.A(n1092), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U1474 (
	.ZN(n1092),
	.B2(\regOut[2][1] ),
	.B1(n936),
	.A2(\regOut[3][1] ),
	.A1(n935), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1475 (
	.ZN(n554),
	.A(\regOut[0][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1476 (
	.ZN(n367),
	.A(\regOut[1][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U1477 (
	.ZN(n1090),
	.C2(n938),
	.C1(n112),
	.B2(n937),
	.B1(n95),
	.A(n1093), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U1478 (
	.ZN(n1093),
	.B2(\regOut[6][1] ),
	.B1(n941),
	.A2(\regOut[7][1] ),
	.A1(n940), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1479 (
	.ZN(n112),
	.A(\regOut[4][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1480 (
	.ZN(n95),
	.A(\regOut[5][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U1481 (
	.ZN(n1089),
	.C2(n943),
	.C1(n44),
	.B2(n942),
	.B1(n20),
	.A(n1094), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U1482 (
	.ZN(n1094),
	.B2(\regOut[10][1] ),
	.B1(n946),
	.A2(\regOut[11][1] ),
	.A1(n945), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1483 (
	.ZN(n44),
	.A(\regOut[8][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1484 (
	.ZN(n20),
	.A(\regOut[9][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U1485 (
	.ZN(n1088),
	.C2(n948),
	.C1(n503),
	.B2(n947),
	.B1(n486),
	.A(n1095), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U1486 (
	.ZN(n1095),
	.B2(\regOut[14][1] ),
	.B1(n951),
	.A2(\regOut[15][1] ),
	.A1(n950), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1487 (
	.ZN(n503),
	.A(\regOut[12][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1488 (
	.ZN(n486),
	.A(\regOut[13][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U1489 (
	.ZN(outA[15]),
	.A2(n1097),
	.A1(n1096), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4_X1 U1490 (
	.ZN(n1097),
	.A4(n1101),
	.A3(n1100),
	.A2(n1099),
	.A1(n1098), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U1491 (
	.ZN(n1101),
	.C2(n909),
	.C1(n436),
	.B2(n908),
	.B1(n419),
	.A(n1102), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U1492 (
	.ZN(n1102),
	.B2(\regOut[18][15] ),
	.B1(n912),
	.A2(\regOut[19][15] ),
	.A1(n911), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1493 (
	.ZN(n436),
	.A(\regOut[16][15] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1494 (
	.ZN(n419),
	.A(\regOut[17][15] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U1495 (
	.ZN(n1100),
	.C2(n914),
	.C1(n351),
	.B2(n913),
	.B1(n334),
	.A(n1103), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U1496 (
	.ZN(n1103),
	.B2(\regOut[22][15] ),
	.B1(n917),
	.A2(\regOut[23][15] ),
	.A1(n916), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1497 (
	.ZN(n351),
	.A(\regOut[20][15] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1498 (
	.ZN(n334),
	.A(\regOut[21][15] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U1499 (
	.ZN(n1099),
	.C2(n919),
	.C1(n283),
	.B2(n918),
	.B1(n266),
	.A(n1104), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U1500 (
	.ZN(n1104),
	.B2(\regOut[26][15] ),
	.B1(n922),
	.A2(\regOut[27][15] ),
	.A1(n921), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1501 (
	.ZN(n283),
	.A(\regOut[24][15] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1502 (
	.ZN(n266),
	.A(\regOut[25][15] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U1503 (
	.ZN(n1098),
	.C2(n924),
	.C1(n164),
	.B2(n923),
	.B1(n147),
	.A(n1105), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U1504 (
	.ZN(n1105),
	.B2(\regOut[28][15] ),
	.B1(n927),
	.A2(\regOut[29][15] ),
	.A1(n926), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1505 (
	.ZN(n164),
	.A(\regOut[30][15] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1506 (
	.ZN(n147),
	.A(\regOut[31][15] ), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4_X1 U1507 (
	.ZN(n1096),
	.A4(n1109),
	.A3(n1108),
	.A2(n1107),
	.A1(n1106), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U1508 (
	.ZN(n1109),
	.C2(n933),
	.C1(n555),
	.B2(n932),
	.B1(n368),
	.A(n1110), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U1509 (
	.ZN(n1110),
	.B2(\regOut[2][15] ),
	.B1(n936),
	.A2(\regOut[3][15] ),
	.A1(n935), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1510 (
	.ZN(n555),
	.A(\regOut[0][15] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1511 (
	.ZN(n368),
	.A(\regOut[1][15] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U1512 (
	.ZN(n1108),
	.C2(n938),
	.C1(n113),
	.B2(n937),
	.B1(n96),
	.A(n1111), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U1513 (
	.ZN(n1111),
	.B2(\regOut[6][15] ),
	.B1(n941),
	.A2(\regOut[7][15] ),
	.A1(n940), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1514 (
	.ZN(n113),
	.A(\regOut[4][15] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1515 (
	.ZN(n96),
	.A(\regOut[5][15] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U1516 (
	.ZN(n1107),
	.C2(n943),
	.C1(n45),
	.B2(n942),
	.B1(n22),
	.A(n1112), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U1517 (
	.ZN(n1112),
	.B2(\regOut[10][15] ),
	.B1(n946),
	.A2(\regOut[11][15] ),
	.A1(n945), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1518 (
	.ZN(n45),
	.A(\regOut[8][15] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1519 (
	.ZN(n22),
	.A(\regOut[9][15] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U1520 (
	.ZN(n1106),
	.C2(n948),
	.C1(n504),
	.B2(n947),
	.B1(n487),
	.A(n1113), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U1521 (
	.ZN(n1113),
	.B2(\regOut[14][15] ),
	.B1(n951),
	.A2(\regOut[15][15] ),
	.A1(n950), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1522 (
	.ZN(n504),
	.A(\regOut[12][15] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1523 (
	.ZN(n487),
	.A(\regOut[13][15] ), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U1524 (
	.ZN(outA[14]),
	.A2(n1115),
	.A1(n1114), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4_X1 U1525 (
	.ZN(n1115),
	.A4(n1119),
	.A3(n1118),
	.A2(n1117),
	.A1(n1116), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U1526 (
	.ZN(n1119),
	.C2(n909),
	.C1(n437),
	.B2(n908),
	.B1(n420),
	.A(n1120), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U1527 (
	.ZN(n1120),
	.B2(\regOut[18][14] ),
	.B1(n912),
	.A2(\regOut[19][14] ),
	.A1(n911), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1528 (
	.ZN(n437),
	.A(\regOut[16][14] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1529 (
	.ZN(n420),
	.A(\regOut[17][14] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U1530 (
	.ZN(n1118),
	.C2(n914),
	.C1(n352),
	.B2(n913),
	.B1(n335),
	.A(n1121), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U1531 (
	.ZN(n1121),
	.B2(\regOut[22][14] ),
	.B1(n917),
	.A2(\regOut[23][14] ),
	.A1(n916), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1532 (
	.ZN(n352),
	.A(\regOut[20][14] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1533 (
	.ZN(n335),
	.A(\regOut[21][14] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U1534 (
	.ZN(n1117),
	.C2(n919),
	.C1(n284),
	.B2(n918),
	.B1(n267),
	.A(n1122), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U1535 (
	.ZN(n1122),
	.B2(\regOut[26][14] ),
	.B1(n922),
	.A2(\regOut[27][14] ),
	.A1(n921), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1536 (
	.ZN(n284),
	.A(\regOut[24][14] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1537 (
	.ZN(n267),
	.A(\regOut[25][14] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U1538 (
	.ZN(n1116),
	.C2(n924),
	.C1(n165),
	.B2(n923),
	.B1(n148),
	.A(n1123), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U1539 (
	.ZN(n1123),
	.B2(\regOut[28][14] ),
	.B1(n927),
	.A2(\regOut[29][14] ),
	.A1(n926), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1540 (
	.ZN(n165),
	.A(\regOut[30][14] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1541 (
	.ZN(n148),
	.A(\regOut[31][14] ), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4_X1 U1542 (
	.ZN(n1114),
	.A4(n1127),
	.A3(n1126),
	.A2(n1125),
	.A1(n1124), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U1543 (
	.ZN(n1127),
	.C2(n933),
	.C1(n556),
	.B2(n932),
	.B1(n369),
	.A(n1128), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U1544 (
	.ZN(n1128),
	.B2(\regOut[2][14] ),
	.B1(n936),
	.A2(\regOut[3][14] ),
	.A1(n935), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1545 (
	.ZN(n556),
	.A(\regOut[0][14] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1546 (
	.ZN(n369),
	.A(\regOut[1][14] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U1547 (
	.ZN(n1126),
	.C2(n938),
	.C1(n114),
	.B2(n937),
	.B1(n97),
	.A(n1129), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U1548 (
	.ZN(n1129),
	.B2(\regOut[6][14] ),
	.B1(n941),
	.A2(\regOut[7][14] ),
	.A1(n940), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1549 (
	.ZN(n114),
	.A(\regOut[4][14] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1550 (
	.ZN(n97),
	.A(\regOut[5][14] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U1551 (
	.ZN(n1125),
	.C2(n943),
	.C1(n46),
	.B2(n942),
	.B1(n24),
	.A(n1130), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U1552 (
	.ZN(n1130),
	.B2(\regOut[10][14] ),
	.B1(n946),
	.A2(\regOut[11][14] ),
	.A1(n945), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1553 (
	.ZN(n46),
	.A(\regOut[8][14] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1554 (
	.ZN(n24),
	.A(\regOut[9][14] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U1555 (
	.ZN(n1124),
	.C2(n948),
	.C1(n505),
	.B2(n947),
	.B1(n488),
	.A(n1131), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U1556 (
	.ZN(n1131),
	.B2(\regOut[14][14] ),
	.B1(n951),
	.A2(\regOut[15][14] ),
	.A1(n950), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1557 (
	.ZN(n505),
	.A(\regOut[12][14] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1558 (
	.ZN(n488),
	.A(\regOut[13][14] ), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U1559 (
	.ZN(outA[13]),
	.A2(n1133),
	.A1(n1132), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4_X1 U1560 (
	.ZN(n1133),
	.A4(n1137),
	.A3(n1136),
	.A2(n1135),
	.A1(n1134), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U1561 (
	.ZN(n1137),
	.C2(n909),
	.C1(n438),
	.B2(n908),
	.B1(n421),
	.A(n1138), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U1562 (
	.ZN(n1138),
	.B2(\regOut[18][13] ),
	.B1(n912),
	.A2(\regOut[19][13] ),
	.A1(n911), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1563 (
	.ZN(n438),
	.A(\regOut[16][13] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1564 (
	.ZN(n421),
	.A(\regOut[17][13] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U1565 (
	.ZN(n1136),
	.C2(n914),
	.C1(n353),
	.B2(n913),
	.B1(n336),
	.A(n1139), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U1566 (
	.ZN(n1139),
	.B2(\regOut[22][13] ),
	.B1(n917),
	.A2(\regOut[23][13] ),
	.A1(n916), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1567 (
	.ZN(n353),
	.A(\regOut[20][13] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1568 (
	.ZN(n336),
	.A(\regOut[21][13] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U1569 (
	.ZN(n1135),
	.C2(n919),
	.C1(n285),
	.B2(n918),
	.B1(n268),
	.A(n1140), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U1570 (
	.ZN(n1140),
	.B2(\regOut[26][13] ),
	.B1(n922),
	.A2(\regOut[27][13] ),
	.A1(n921), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1571 (
	.ZN(n285),
	.A(\regOut[24][13] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1572 (
	.ZN(n268),
	.A(\regOut[25][13] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U1573 (
	.ZN(n1134),
	.C2(n924),
	.C1(n166),
	.B2(n923),
	.B1(n149),
	.A(n1141), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U1574 (
	.ZN(n1141),
	.B2(\regOut[28][13] ),
	.B1(n927),
	.A2(\regOut[29][13] ),
	.A1(n926), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1575 (
	.ZN(n166),
	.A(\regOut[30][13] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1576 (
	.ZN(n149),
	.A(\regOut[31][13] ), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4_X1 U1577 (
	.ZN(n1132),
	.A4(n1145),
	.A3(n1144),
	.A2(n1143),
	.A1(n1142), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U1578 (
	.ZN(n1145),
	.C2(n933),
	.C1(n557),
	.B2(n932),
	.B1(n370),
	.A(n1146), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U1579 (
	.ZN(n1146),
	.B2(\regOut[2][13] ),
	.B1(n936),
	.A2(\regOut[3][13] ),
	.A1(n935), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1580 (
	.ZN(n557),
	.A(\regOut[0][13] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1581 (
	.ZN(n370),
	.A(\regOut[1][13] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U1582 (
	.ZN(n1144),
	.C2(n938),
	.C1(n115),
	.B2(n937),
	.B1(n98),
	.A(n1147), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U1583 (
	.ZN(n1147),
	.B2(\regOut[6][13] ),
	.B1(n941),
	.A2(\regOut[7][13] ),
	.A1(n940), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1584 (
	.ZN(n115),
	.A(\regOut[4][13] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1585 (
	.ZN(n98),
	.A(\regOut[5][13] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U1586 (
	.ZN(n1143),
	.C2(n943),
	.C1(n47),
	.B2(n942),
	.B1(n26),
	.A(n1148), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U1587 (
	.ZN(n1148),
	.B2(\regOut[10][13] ),
	.B1(n946),
	.A2(\regOut[11][13] ),
	.A1(n945), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1588 (
	.ZN(n47),
	.A(\regOut[8][13] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1589 (
	.ZN(n26),
	.A(\regOut[9][13] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U1590 (
	.ZN(n1142),
	.C2(n948),
	.C1(n506),
	.B2(n947),
	.B1(n489),
	.A(n1149), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U1591 (
	.ZN(n1149),
	.B2(\regOut[14][13] ),
	.B1(n951),
	.A2(\regOut[15][13] ),
	.A1(n950), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1592 (
	.ZN(n506),
	.A(\regOut[12][13] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1593 (
	.ZN(n489),
	.A(\regOut[13][13] ), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U1594 (
	.ZN(outA[12]),
	.A2(n1151),
	.A1(n1150), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4_X1 U1595 (
	.ZN(n1151),
	.A4(n1155),
	.A3(n1154),
	.A2(n1153),
	.A1(n1152), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U1596 (
	.ZN(n1155),
	.C2(n909),
	.C1(n439),
	.B2(n908),
	.B1(n422),
	.A(n1156), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U1597 (
	.ZN(n1156),
	.B2(\regOut[18][12] ),
	.B1(n912),
	.A2(\regOut[19][12] ),
	.A1(n911), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1598 (
	.ZN(n439),
	.A(\regOut[16][12] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1599 (
	.ZN(n422),
	.A(\regOut[17][12] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U1600 (
	.ZN(n1154),
	.C2(n914),
	.C1(n354),
	.B2(n913),
	.B1(n337),
	.A(n1157), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U1601 (
	.ZN(n1157),
	.B2(\regOut[22][12] ),
	.B1(n917),
	.A2(\regOut[23][12] ),
	.A1(n916), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1602 (
	.ZN(n354),
	.A(\regOut[20][12] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1603 (
	.ZN(n337),
	.A(\regOut[21][12] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U1604 (
	.ZN(n1153),
	.C2(n919),
	.C1(n286),
	.B2(n918),
	.B1(n269),
	.A(n1158), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U1605 (
	.ZN(n1158),
	.B2(\regOut[26][12] ),
	.B1(n922),
	.A2(\regOut[27][12] ),
	.A1(n921), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1606 (
	.ZN(n286),
	.A(\regOut[24][12] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1607 (
	.ZN(n269),
	.A(\regOut[25][12] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U1608 (
	.ZN(n1152),
	.C2(n924),
	.C1(n167),
	.B2(n923),
	.B1(n150),
	.A(n1159), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U1609 (
	.ZN(n1159),
	.B2(\regOut[28][12] ),
	.B1(n927),
	.A2(\regOut[29][12] ),
	.A1(n926), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1610 (
	.ZN(n167),
	.A(\regOut[30][12] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1611 (
	.ZN(n150),
	.A(\regOut[31][12] ), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4_X1 U1612 (
	.ZN(n1150),
	.A4(n1163),
	.A3(n1162),
	.A2(n1161),
	.A1(n1160), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U1613 (
	.ZN(n1163),
	.C2(n933),
	.C1(n558),
	.B2(n932),
	.B1(n371),
	.A(n1164), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U1614 (
	.ZN(n1164),
	.B2(\regOut[2][12] ),
	.B1(n936),
	.A2(\regOut[3][12] ),
	.A1(n935), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1615 (
	.ZN(n558),
	.A(\regOut[0][12] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1616 (
	.ZN(n371),
	.A(\regOut[1][12] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U1617 (
	.ZN(n1162),
	.C2(n938),
	.C1(n116),
	.B2(n937),
	.B1(n99),
	.A(n1165), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U1618 (
	.ZN(n1165),
	.B2(\regOut[6][12] ),
	.B1(n941),
	.A2(\regOut[7][12] ),
	.A1(n940), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1619 (
	.ZN(n116),
	.A(\regOut[4][12] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1620 (
	.ZN(n99),
	.A(\regOut[5][12] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U1621 (
	.ZN(n1161),
	.C2(n943),
	.C1(n48),
	.B2(n942),
	.B1(n28),
	.A(n1166), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U1622 (
	.ZN(n1166),
	.B2(\regOut[10][12] ),
	.B1(n946),
	.A2(\regOut[11][12] ),
	.A1(n945), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1623 (
	.ZN(n48),
	.A(\regOut[8][12] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1624 (
	.ZN(n28),
	.A(\regOut[9][12] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U1625 (
	.ZN(n1160),
	.C2(n948),
	.C1(n507),
	.B2(n947),
	.B1(n490),
	.A(n1167), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U1626 (
	.ZN(n1167),
	.B2(\regOut[14][12] ),
	.B1(n951),
	.A2(\regOut[15][12] ),
	.A1(n950), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1627 (
	.ZN(n507),
	.A(\regOut[12][12] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1628 (
	.ZN(n490),
	.A(\regOut[13][12] ), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U1629 (
	.ZN(outA[11]),
	.A2(n1169),
	.A1(n1168), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4_X1 U1630 (
	.ZN(n1169),
	.A4(n1173),
	.A3(n1172),
	.A2(n1171),
	.A1(n1170), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U1631 (
	.ZN(n1173),
	.C2(n909),
	.C1(n440),
	.B2(n908),
	.B1(n423),
	.A(n1174), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U1632 (
	.ZN(n1174),
	.B2(\regOut[18][11] ),
	.B1(n912),
	.A2(\regOut[19][11] ),
	.A1(n911), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1633 (
	.ZN(n440),
	.A(\regOut[16][11] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1634 (
	.ZN(n423),
	.A(\regOut[17][11] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U1635 (
	.ZN(n1172),
	.C2(n914),
	.C1(n355),
	.B2(n913),
	.B1(n338),
	.A(n1175), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U1636 (
	.ZN(n1175),
	.B2(\regOut[22][11] ),
	.B1(n917),
	.A2(\regOut[23][11] ),
	.A1(n916), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1637 (
	.ZN(n355),
	.A(\regOut[20][11] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1638 (
	.ZN(n338),
	.A(\regOut[21][11] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U1639 (
	.ZN(n1171),
	.C2(n919),
	.C1(n287),
	.B2(n918),
	.B1(n270),
	.A(n1176), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U1640 (
	.ZN(n1176),
	.B2(\regOut[26][11] ),
	.B1(n922),
	.A2(\regOut[27][11] ),
	.A1(n921), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1641 (
	.ZN(n287),
	.A(\regOut[24][11] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1642 (
	.ZN(n270),
	.A(\regOut[25][11] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U1643 (
	.ZN(n1170),
	.C2(n924),
	.C1(n168),
	.B2(n923),
	.B1(n151),
	.A(n1177), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U1644 (
	.ZN(n1177),
	.B2(\regOut[28][11] ),
	.B1(n927),
	.A2(\regOut[29][11] ),
	.A1(n926), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1645 (
	.ZN(n168),
	.A(\regOut[30][11] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1646 (
	.ZN(n151),
	.A(\regOut[31][11] ), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4_X1 U1647 (
	.ZN(n1168),
	.A4(n1181),
	.A3(n1180),
	.A2(n1179),
	.A1(n1178), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U1648 (
	.ZN(n1181),
	.C2(n933),
	.C1(n559),
	.B2(n932),
	.B1(n372),
	.A(n1182), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U1649 (
	.ZN(n1182),
	.B2(\regOut[2][11] ),
	.B1(n936),
	.A2(\regOut[3][11] ),
	.A1(n935), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1650 (
	.ZN(n559),
	.A(\regOut[0][11] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1651 (
	.ZN(n372),
	.A(\regOut[1][11] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U1652 (
	.ZN(n1180),
	.C2(n938),
	.C1(n117),
	.B2(n937),
	.B1(n100),
	.A(n1183), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U1653 (
	.ZN(n1183),
	.B2(\regOut[6][11] ),
	.B1(n941),
	.A2(\regOut[7][11] ),
	.A1(n940), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1654 (
	.ZN(n117),
	.A(\regOut[4][11] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1655 (
	.ZN(n100),
	.A(\regOut[5][11] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U1656 (
	.ZN(n1179),
	.C2(n943),
	.C1(n49),
	.B2(n942),
	.B1(n30),
	.A(n1184), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U1657 (
	.ZN(n1184),
	.B2(\regOut[10][11] ),
	.B1(n946),
	.A2(\regOut[11][11] ),
	.A1(n945), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1658 (
	.ZN(n49),
	.A(\regOut[8][11] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1659 (
	.ZN(n30),
	.A(\regOut[9][11] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U1660 (
	.ZN(n1178),
	.C2(n948),
	.C1(n508),
	.B2(n947),
	.B1(n491),
	.A(n1185), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U1661 (
	.ZN(n1185),
	.B2(\regOut[14][11] ),
	.B1(n951),
	.A2(\regOut[15][11] ),
	.A1(n950), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1662 (
	.ZN(n508),
	.A(\regOut[12][11] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1663 (
	.ZN(n491),
	.A(\regOut[13][11] ), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U1664 (
	.ZN(outA[10]),
	.A2(n1187),
	.A1(n1186), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4_X1 U1665 (
	.ZN(n1187),
	.A4(n1191),
	.A3(n1190),
	.A2(n1189),
	.A1(n1188), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U1666 (
	.ZN(n1191),
	.C2(n909),
	.C1(n441),
	.B2(n908),
	.B1(n424),
	.A(n1192), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U1667 (
	.ZN(n1192),
	.B2(\regOut[18][10] ),
	.B1(n912),
	.A2(\regOut[19][10] ),
	.A1(n911), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1668 (
	.ZN(n441),
	.A(\regOut[16][10] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1669 (
	.ZN(n424),
	.A(\regOut[17][10] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U1670 (
	.ZN(n1190),
	.C2(n914),
	.C1(n356),
	.B2(n913),
	.B1(n339),
	.A(n1193), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U1671 (
	.ZN(n1193),
	.B2(\regOut[22][10] ),
	.B1(n917),
	.A2(\regOut[23][10] ),
	.A1(n916), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1672 (
	.ZN(n356),
	.A(\regOut[20][10] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1673 (
	.ZN(n339),
	.A(\regOut[21][10] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U1674 (
	.ZN(n1189),
	.C2(n919),
	.C1(n288),
	.B2(n918),
	.B1(n271),
	.A(n1194), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U1675 (
	.ZN(n1194),
	.B2(\regOut[26][10] ),
	.B1(n922),
	.A2(\regOut[27][10] ),
	.A1(n921), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1676 (
	.ZN(n288),
	.A(\regOut[24][10] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1677 (
	.ZN(n271),
	.A(\regOut[25][10] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U1678 (
	.ZN(n1188),
	.C2(n924),
	.C1(n169),
	.B2(n923),
	.B1(n152),
	.A(n1195), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U1679 (
	.ZN(n1195),
	.B2(\regOut[28][10] ),
	.B1(n927),
	.A2(\regOut[29][10] ),
	.A1(n926), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1680 (
	.ZN(n169),
	.A(\regOut[30][10] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1681 (
	.ZN(n152),
	.A(\regOut[31][10] ), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4_X1 U1682 (
	.ZN(n1186),
	.A4(n1199),
	.A3(n1198),
	.A2(n1197),
	.A1(n1196), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U1683 (
	.ZN(n1199),
	.C2(n933),
	.C1(n560),
	.B2(n932),
	.B1(n373),
	.A(n1200), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U1684 (
	.ZN(n1200),
	.B2(\regOut[2][10] ),
	.B1(n936),
	.A2(\regOut[3][10] ),
	.A1(n935), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1685 (
	.ZN(n560),
	.A(\regOut[0][10] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1686 (
	.ZN(n373),
	.A(\regOut[1][10] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U1687 (
	.ZN(n1198),
	.C2(n938),
	.C1(n118),
	.B2(n937),
	.B1(n101),
	.A(n1201), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U1688 (
	.ZN(n1201),
	.B2(\regOut[6][10] ),
	.B1(n941),
	.A2(\regOut[7][10] ),
	.A1(n940), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1689 (
	.ZN(n118),
	.A(\regOut[4][10] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1690 (
	.ZN(n101),
	.A(\regOut[5][10] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U1691 (
	.ZN(n1197),
	.C2(n943),
	.C1(n50),
	.B2(n942),
	.B1(n32),
	.A(n1202), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U1692 (
	.ZN(n1202),
	.B2(\regOut[10][10] ),
	.B1(n946),
	.A2(\regOut[11][10] ),
	.A1(n945), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1693 (
	.ZN(n50),
	.A(\regOut[8][10] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1694 (
	.ZN(n32),
	.A(\regOut[9][10] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U1695 (
	.ZN(n1196),
	.C2(n948),
	.C1(n509),
	.B2(n947),
	.B1(n492),
	.A(n1203), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U1696 (
	.ZN(n1203),
	.B2(\regOut[14][10] ),
	.B1(n951),
	.A2(\regOut[15][10] ),
	.A1(n950), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1697 (
	.ZN(n509),
	.A(\regOut[12][10] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1698 (
	.ZN(n492),
	.A(\regOut[13][10] ), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U1699 (
	.ZN(outA[0]),
	.A2(n1205),
	.A1(n1204), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4_X1 U1700 (
	.ZN(n1205),
	.A4(n1209),
	.A3(n1208),
	.A2(n1207),
	.A1(n1206), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U1701 (
	.ZN(n1209),
	.C2(n909),
	.C1(n442),
	.B2(n908),
	.B1(n425),
	.A(n1210), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U1702 (
	.ZN(n1210),
	.B2(\regOut[18][0] ),
	.B1(n912),
	.A2(\regOut[19][0] ),
	.A1(n911), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2_X1 U1703 (
	.ZN(n912),
	.A2(n1212),
	.A1(n1211), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2_X1 U1704 (
	.ZN(n911),
	.A2(n1212),
	.A1(n1213), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U1705 (
	.ZN(n909),
	.A2(n1214),
	.A1(n1211), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1706 (
	.ZN(n442),
	.A(\regOut[16][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U1707 (
	.ZN(n908),
	.A2(n1214),
	.A1(n1213), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1708 (
	.ZN(n425),
	.A(\regOut[17][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U1709 (
	.ZN(n1208),
	.C2(n914),
	.C1(n357),
	.B2(n913),
	.B1(n340),
	.A(n1215), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U1710 (
	.ZN(n1215),
	.B2(\regOut[22][0] ),
	.B1(n917),
	.A2(\regOut[23][0] ),
	.A1(n916), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2_X1 U1711 (
	.ZN(n917),
	.A2(n1216),
	.A1(n1211), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2_X1 U1712 (
	.ZN(n916),
	.A2(n1216),
	.A1(n1213), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U1713 (
	.ZN(n914),
	.A2(n1217),
	.A1(n1211), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2_X1 U1714 (
	.ZN(n1211),
	.A2(n1219),
	.A1(n1218), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1715 (
	.ZN(n357),
	.A(\regOut[20][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U1716 (
	.ZN(n913),
	.A2(n1217),
	.A1(n1213), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2_X1 U1717 (
	.ZN(n1213),
	.A2(addressA[0]),
	.A1(n1218), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2_X1 U1718 (
	.ZN(n1218),
	.A2(n1220),
	.A1(addressA[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1719 (
	.ZN(n340),
	.A(\regOut[21][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U1720 (
	.ZN(n1207),
	.C2(n919),
	.C1(n289),
	.B2(n918),
	.B1(n272),
	.A(n1221), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U1721 (
	.ZN(n1221),
	.B2(\regOut[26][0] ),
	.B1(n922),
	.A2(\regOut[27][0] ),
	.A1(n921), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2_X1 U1722 (
	.ZN(n922),
	.A2(n1222),
	.A1(n1212), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2_X1 U1723 (
	.ZN(n921),
	.A2(n1223),
	.A1(n1212), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U1724 (
	.ZN(n919),
	.A2(n1222),
	.A1(n1214), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1725 (
	.ZN(n289),
	.A(\regOut[24][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U1726 (
	.ZN(n918),
	.A2(n1223),
	.A1(n1214), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1727 (
	.ZN(n272),
	.A(\regOut[25][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U1728 (
	.ZN(n1206),
	.C2(n924),
	.C1(n170),
	.B2(n923),
	.B1(n153),
	.A(n1224), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U1729 (
	.ZN(n1224),
	.B2(\regOut[28][0] ),
	.B1(n927),
	.A2(\regOut[29][0] ),
	.A1(n926), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2_X1 U1730 (
	.ZN(n927),
	.A2(n1222),
	.A1(n1217), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2_X1 U1731 (
	.ZN(n926),
	.A2(n1223),
	.A1(n1217), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U1732 (
	.ZN(n924),
	.A2(n1216),
	.A1(n1222), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2_X1 U1733 (
	.ZN(n1222),
	.A2(n1219),
	.A1(n1225), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1734 (
	.ZN(n170),
	.A(\regOut[30][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U1735 (
	.ZN(n923),
	.A2(n1223),
	.A1(n1216), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2_X1 U1736 (
	.ZN(n1223),
	.A2(n1225),
	.A1(addressA[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2_X1 U1737 (
	.ZN(n1225),
	.A2(addressA[3]),
	.A1(addressA[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1738 (
	.ZN(n153),
	.A(\regOut[31][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4_X1 U1739 (
	.ZN(n1204),
	.A4(n1229),
	.A3(n1228),
	.A2(n1227),
	.A1(n1226), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U1740 (
	.ZN(n1229),
	.C2(n933),
	.C1(n561),
	.B2(n932),
	.B1(n374),
	.A(n1230), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U1741 (
	.ZN(n1230),
	.B2(\regOut[2][0] ),
	.B1(n936),
	.A2(\regOut[3][0] ),
	.A1(n935), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2_X1 U1742 (
	.ZN(n936),
	.A2(n1212),
	.A1(n1231), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2_X1 U1743 (
	.ZN(n935),
	.A2(n1212),
	.A1(n1232), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U1744 (
	.ZN(n933),
	.A2(n1214),
	.A1(n1231), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1745 (
	.ZN(n561),
	.A(\regOut[0][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U1746 (
	.ZN(n932),
	.A2(n1214),
	.A1(n1232), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1747 (
	.ZN(n374),
	.A(\regOut[1][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U1748 (
	.ZN(n1228),
	.C2(n938),
	.C1(n119),
	.B2(n937),
	.B1(n102),
	.A(n1233), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U1749 (
	.ZN(n1233),
	.B2(\regOut[6][0] ),
	.B1(n941),
	.A2(\regOut[7][0] ),
	.A1(n940), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2_X1 U1750 (
	.ZN(n941),
	.A2(n1216),
	.A1(n1231), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2_X1 U1751 (
	.ZN(n940),
	.A2(n1216),
	.A1(n1232), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U1752 (
	.ZN(n938),
	.A2(n1217),
	.A1(n1231), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2_X1 U1753 (
	.ZN(n1231),
	.A2(n1219),
	.A1(n1234), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1754 (
	.ZN(n119),
	.A(\regOut[4][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U1755 (
	.ZN(n937),
	.A2(n1217),
	.A1(n1232), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2_X1 U1756 (
	.ZN(n1232),
	.A2(addressA[0]),
	.A1(n1234), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2_X1 U1757 (
	.ZN(n1234),
	.A2(addressA[4]),
	.A1(addressA[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1758 (
	.ZN(n102),
	.A(\regOut[5][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U1759 (
	.ZN(n1227),
	.C2(n943),
	.C1(n51),
	.B2(n942),
	.B1(n34),
	.A(n1235), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U1760 (
	.ZN(n1235),
	.B2(\regOut[10][0] ),
	.B1(n946),
	.A2(\regOut[11][0] ),
	.A1(n945), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2_X1 U1761 (
	.ZN(n946),
	.A2(n1212),
	.A1(n1236), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2_X1 U1762 (
	.ZN(n945),
	.A2(n1212),
	.A1(n1237), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2_X1 U1763 (
	.ZN(n1212),
	.A2(addressA[2]),
	.A1(n1238), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U1764 (
	.ZN(n943),
	.A2(n1214),
	.A1(n1236), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1765 (
	.ZN(n51),
	.A(\regOut[8][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U1766 (
	.ZN(n942),
	.A2(n1214),
	.A1(n1237), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2_X2 U1767 (
	.ZN(n1214),
	.A2(addressA[2]),
	.A1(addressA[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1768 (
	.ZN(n34),
	.A(\regOut[9][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221_X1 U1769 (
	.ZN(n1226),
	.C2(n948),
	.C1(n510),
	.B2(n947),
	.B1(n493),
	.A(n1239), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22_X1 U1770 (
	.ZN(n1239),
	.B2(\regOut[14][0] ),
	.B1(n951),
	.A2(\regOut[15][0] ),
	.A1(n950), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2_X1 U1771 (
	.ZN(n951),
	.A2(n1216),
	.A1(n1236), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2_X1 U1772 (
	.ZN(n950),
	.A2(n1216),
	.A1(n1237), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2_X1 U1773 (
	.ZN(n1216),
	.A2(n1238),
	.A1(n1240), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1774 (
	.ZN(n1238),
	.A(addressA[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U1775 (
	.ZN(n948),
	.A2(n1217),
	.A1(n1236), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2_X1 U1776 (
	.ZN(n1236),
	.A2(n1219),
	.A1(n1241), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1777 (
	.ZN(n1219),
	.A(addressA[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1778 (
	.ZN(n510),
	.A(\regOut[12][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2_X1 U1779 (
	.ZN(n947),
	.A2(n1217),
	.A1(n1237), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2_X2 U1780 (
	.ZN(n1217),
	.A2(addressA[1]),
	.A1(n1240), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1781 (
	.ZN(n1240),
	.A(addressA[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2_X1 U1782 (
	.ZN(n1237),
	.A2(addressA[0]),
	.A1(n1241), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2_X1 U1783 (
	.ZN(n1241),
	.A2(addressA[4]),
	.A1(n1220), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1784 (
	.ZN(n1220),
	.A(addressA[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1785 (
	.ZN(n493),
	.A(\regOut[13][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   SingleReg_31 RegX_0 (
	.data({ \regIn[0][15] ,
		\regIn[0][14] ,
		\regIn[0][13] ,
		\regIn[0][12] ,
		\regIn[0][11] ,
		\regIn[0][10] ,
		\regIn[0][9] ,
		\regIn[0][8] ,
		\regIn[0][7] ,
		\regIn[0][6] ,
		\regIn[0][5] ,
		\regIn[0][4] ,
		\regIn[0][3] ,
		\regIn[0][2] ,
		\regIn[0][1] ,
		\regIn[0][0]  }),
	.clk(clk__L2_N2),
	.reset(reset),
	.write(write),
	.dataOut({ \regOut[0][15] ,
		\regOut[0][14] ,
		\regOut[0][13] ,
		\regOut[0][12] ,
		\regOut[0][11] ,
		\regOut[0][10] ,
		\regOut[0][9] ,
		\regOut[0][8] ,
		\regOut[0][7] ,
		\regOut[0][6] ,
		\regOut[0][5] ,
		\regOut[0][4] ,
		\regOut[0][3] ,
		\regOut[0][2] ,
		\regOut[0][1] ,
		\regOut[0][0]  }),
	.FE_OFN1_write(FE_OFN21_write),
	.FE_OFN2_write(FE_OFN41_write),
	.FE_OFN18_write(FE_OFN18_write),
	.FE_OFN20_write(FE_OFN20_write),
	.FE_OFN22_write(FE_OFN22_write),
	.FE_OFN24_write(FE_OFN24_write),
	.FE_OFN29_write(FE_OFN29_write),
	.FE_OFN31_write(FE_OFN31_write),
	.clk__L2_N3(clk__L2_N3),
	.clk__L2_N4(clk__L2_N4),
	.clk__L2_N7(clk__L2_N7),
	.clk__L2_N8(clk__L2_N8), 
	.VDD(VDD), 
	.VSS(VSS));
   SingleReg_30 RegX_1 (
	.data({ \regIn[1][15] ,
		\regIn[1][14] ,
		\regIn[1][13] ,
		\regIn[1][12] ,
		\regIn[1][11] ,
		\regIn[1][10] ,
		\regIn[1][9] ,
		\regIn[1][8] ,
		\regIn[1][7] ,
		\regIn[1][6] ,
		\regIn[1][5] ,
		\regIn[1][4] ,
		\regIn[1][3] ,
		\regIn[1][2] ,
		\regIn[1][1] ,
		\regIn[1][0]  }),
	.clk(clk__L2_N2),
	.reset(reset),
	.write(write),
	.dataOut({ \regOut[1][15] ,
		\regOut[1][14] ,
		\regOut[1][13] ,
		\regOut[1][12] ,
		\regOut[1][11] ,
		\regOut[1][10] ,
		\regOut[1][9] ,
		\regOut[1][8] ,
		\regOut[1][7] ,
		\regOut[1][6] ,
		\regOut[1][5] ,
		\regOut[1][4] ,
		\regOut[1][3] ,
		\regOut[1][2] ,
		\regOut[1][1] ,
		\regOut[1][0]  }),
	.FE_OFN1_write(write),
	.FE_OFN2_write(FE_OFN41_write),
	.FE_OFN18_write(FE_OFN18_write),
	.FE_OFN20_write(FE_OFN20_write),
	.FE_OFN22_write(FE_OFN22_write),
	.FE_OFN29_write(FE_OFN29_write),
	.FE_OFN31_write(FE_OFN31_write),
	.clk__L2_N3(clk__L2_N3),
	.clk__L2_N4(clk__L2_N4),
	.clk__L2_N7(clk__L2_N7),
	.clk__L2_N8(clk__L2_N8), 
	.VDD(VDD), 
	.VSS(VSS));
   SingleReg_29 RegX_2 (
	.data({ \regIn[2][15] ,
		\regIn[2][14] ,
		\regIn[2][13] ,
		\regIn[2][12] ,
		\regIn[2][11] ,
		\regIn[2][10] ,
		\regIn[2][9] ,
		\regIn[2][8] ,
		\regIn[2][7] ,
		\regIn[2][6] ,
		\regIn[2][5] ,
		\regIn[2][4] ,
		\regIn[2][3] ,
		\regIn[2][2] ,
		\regIn[2][1] ,
		\regIn[2][0]  }),
	.clk(clk__L2_N7),
	.reset(reset),
	.write(write),
	.dataOut({ \regOut[2][15] ,
		\regOut[2][14] ,
		\regOut[2][13] ,
		\regOut[2][12] ,
		\regOut[2][11] ,
		\regOut[2][10] ,
		\regOut[2][9] ,
		\regOut[2][8] ,
		\regOut[2][7] ,
		\regOut[2][6] ,
		\regOut[2][5] ,
		\regOut[2][4] ,
		\regOut[2][3] ,
		\regOut[2][2] ,
		\regOut[2][1] ,
		\regOut[2][0]  }),
	.FE_OFN0_write(write),
	.FE_OFN15_write(FE_OFN15_write),
	.FE_OFN16_write(FE_OFN16_write),
	.FE_OFN17_write(FE_OFN17_write),
	.clk__L2_N8(clk__L2_N8), 
	.VDD(VDD), 
	.VSS(VSS));
   SingleReg_28 RegX_3 (
	.data({ \regIn[3][15] ,
		\regIn[3][14] ,
		\regIn[3][13] ,
		\regIn[3][12] ,
		\regIn[3][11] ,
		\regIn[3][10] ,
		\regIn[3][9] ,
		\regIn[3][8] ,
		\regIn[3][7] ,
		\regIn[3][6] ,
		\regIn[3][5] ,
		\regIn[3][4] ,
		\regIn[3][3] ,
		\regIn[3][2] ,
		\regIn[3][1] ,
		\regIn[3][0]  }),
	.clk(clk__L2_N7),
	.reset(reset),
	.write(FE_OFN16_write),
	.dataOut({ \regOut[3][15] ,
		\regOut[3][14] ,
		\regOut[3][13] ,
		\regOut[3][12] ,
		\regOut[3][11] ,
		\regOut[3][10] ,
		\regOut[3][9] ,
		\regOut[3][8] ,
		\regOut[3][7] ,
		\regOut[3][6] ,
		\regOut[3][5] ,
		\regOut[3][4] ,
		\regOut[3][3] ,
		\regOut[3][2] ,
		\regOut[3][1] ,
		\regOut[3][0]  }),
	.FE_OFN0_write(write),
	.FE_OFN17_write(FE_OFN17_write),
	.FE_OFN18_write(FE_OFN18_write),
	.FE_OFN20_write(FE_OFN20_write),
	.clk__L2_N8(clk__L2_N8), 
	.VDD(VDD), 
	.VSS(VSS));
   SingleReg_27 RegX_4 (
	.data({ \regIn[4][15] ,
		\regIn[4][14] ,
		\regIn[4][13] ,
		\regIn[4][12] ,
		\regIn[4][11] ,
		\regIn[4][10] ,
		\regIn[4][9] ,
		\regIn[4][8] ,
		\regIn[4][7] ,
		\regIn[4][6] ,
		\regIn[4][5] ,
		\regIn[4][4] ,
		\regIn[4][3] ,
		\regIn[4][2] ,
		\regIn[4][1] ,
		\regIn[4][0]  }),
	.clk(clk__L2_N0),
	.reset(reset),
	.write(FE_OFN21_write),
	.dataOut({ \regOut[4][15] ,
		\regOut[4][14] ,
		\regOut[4][13] ,
		\regOut[4][12] ,
		\regOut[4][11] ,
		\regOut[4][10] ,
		\regOut[4][9] ,
		\regOut[4][8] ,
		\regOut[4][7] ,
		\regOut[4][6] ,
		\regOut[4][5] ,
		\regOut[4][4] ,
		\regOut[4][3] ,
		\regOut[4][2] ,
		\regOut[4][1] ,
		\regOut[4][0]  }),
	.FE_OFN5_write(FE_OFN49_write),
	.FE_OFN6_write(FE_OFN32_write),
	.FE_OFN32_write(FE_OFN32_write),
	.FE_OFN36_write(FE_UNCONNECTED_0),
	.FE_OFN44_write(FE_OFN44_write),
	.clk__L2_N2(clk__L2_N2),
	.clk__L2_N3(clk__L2_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   SingleReg_26 RegX_5 (
	.data({ \regIn[5][15] ,
		\regIn[5][14] ,
		\regIn[5][13] ,
		\regIn[5][12] ,
		\regIn[5][11] ,
		\regIn[5][10] ,
		\regIn[5][9] ,
		\regIn[5][8] ,
		\regIn[5][7] ,
		\regIn[5][6] ,
		\regIn[5][5] ,
		\regIn[5][4] ,
		\regIn[5][3] ,
		\regIn[5][2] ,
		\regIn[5][1] ,
		\regIn[5][0]  }),
	.clk(clk__L2_N0),
	.reset(reset),
	.write(FE_OFN21_write),
	.dataOut({ \regOut[5][15] ,
		\regOut[5][14] ,
		\regOut[5][13] ,
		\regOut[5][12] ,
		\regOut[5][11] ,
		\regOut[5][10] ,
		\regOut[5][9] ,
		\regOut[5][8] ,
		\regOut[5][7] ,
		\regOut[5][6] ,
		\regOut[5][5] ,
		\regOut[5][4] ,
		\regOut[5][3] ,
		\regOut[5][2] ,
		\regOut[5][1] ,
		\regOut[5][0]  }),
	.FE_OFN5_write(FE_OFN49_write),
	.FE_OFN6_write(FE_OFN44_write),
	.FE_OFN32_write(FE_OFN32_write),
	.FE_OFN36_write(FE_UNCONNECTED_0),
	.clk__L2_N2(clk__L2_N2),
	.clk__L2_N3(clk__L2_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   SingleReg_25 RegX_6 (
	.data({ \regIn[6][15] ,
		\regIn[6][14] ,
		\regIn[6][13] ,
		\regIn[6][12] ,
		\regIn[6][11] ,
		\regIn[6][10] ,
		\regIn[6][9] ,
		\regIn[6][8] ,
		\regIn[6][7] ,
		\regIn[6][6] ,
		\regIn[6][5] ,
		\regIn[6][4] ,
		\regIn[6][3] ,
		\regIn[6][2] ,
		\regIn[6][1] ,
		\regIn[6][0]  }),
	.clk(clk__L2_N0),
	.reset(reset),
	.write(FE_OFN21_write),
	.dataOut({ \regOut[6][15] ,
		\regOut[6][14] ,
		\regOut[6][13] ,
		\regOut[6][12] ,
		\regOut[6][11] ,
		\regOut[6][10] ,
		\regOut[6][9] ,
		\regOut[6][8] ,
		\regOut[6][7] ,
		\regOut[6][6] ,
		\regOut[6][5] ,
		\regOut[6][4] ,
		\regOut[6][3] ,
		\regOut[6][2] ,
		\regOut[6][1] ,
		\regOut[6][0]  }),
	.FE_OFN2_write(FE_OFN21_write),
	.FE_OFN6_write(FE_OFN32_write),
	.FE_OFN25_write(FE_OFN25_write),
	.FE_OFN31_write(FE_OFN31_write),
	.FE_OFN32_write(FE_OFN32_write),
	.FE_OFN41_write(FE_OFN41_write),
	.clk__L2_N2(clk__L2_N2),
	.clk__L2_N3(clk__L2_N3),
	.clk__L2_N4(clk__L2_N4), 
	.VDD(VDD), 
	.VSS(VSS));
   SingleReg_24 RegX_7 (
	.data({ \regIn[7][15] ,
		\regIn[7][14] ,
		\regIn[7][13] ,
		\regIn[7][12] ,
		\regIn[7][11] ,
		\regIn[7][10] ,
		\regIn[7][9] ,
		\regIn[7][8] ,
		\regIn[7][7] ,
		\regIn[7][6] ,
		\regIn[7][5] ,
		\regIn[7][4] ,
		\regIn[7][3] ,
		\regIn[7][2] ,
		\regIn[7][1] ,
		\regIn[7][0]  }),
	.clk(clk__L2_N0),
	.reset(reset),
	.write(FE_OFN21_write),
	.dataOut({ \regOut[7][15] ,
		\regOut[7][14] ,
		\regOut[7][13] ,
		\regOut[7][12] ,
		\regOut[7][11] ,
		\regOut[7][10] ,
		\regOut[7][9] ,
		\regOut[7][8] ,
		\regOut[7][7] ,
		\regOut[7][6] ,
		\regOut[7][5] ,
		\regOut[7][4] ,
		\regOut[7][3] ,
		\regOut[7][2] ,
		\regOut[7][1] ,
		\regOut[7][0]  }),
	.FE_OFN2_write(FE_OFN41_write),
	.FE_OFN24_write(FE_OFN24_write),
	.FE_OFN25_write(FE_OFN25_write),
	.FE_OFN31_write(FE_OFN31_write),
	.clk__L2_N2(clk__L2_N2),
	.clk__L2_N3(clk__L2_N3),
	.clk__L2_N4(clk__L2_N4), 
	.VDD(VDD), 
	.VSS(VSS));
   SingleReg_23 RegX_8 (
	.data({ \regIn[8][15] ,
		\regIn[8][14] ,
		\regIn[8][13] ,
		\regIn[8][12] ,
		\regIn[8][11] ,
		\regIn[8][10] ,
		\regIn[8][9] ,
		\regIn[8][8] ,
		\regIn[8][7] ,
		\regIn[8][6] ,
		\regIn[8][5] ,
		\regIn[8][4] ,
		\regIn[8][3] ,
		\regIn[8][2] ,
		\regIn[8][1] ,
		\regIn[8][0]  }),
	.clk(clk__L2_N0),
	.reset(reset),
	.write(FE_OFN32_write),
	.dataOut({ \regOut[8][15] ,
		\regOut[8][14] ,
		\regOut[8][13] ,
		\regOut[8][12] ,
		\regOut[8][11] ,
		\regOut[8][10] ,
		\regOut[8][9] ,
		\regOut[8][8] ,
		\regOut[8][7] ,
		\regOut[8][6] ,
		\regOut[8][5] ,
		\regOut[8][4] ,
		\regOut[8][3] ,
		\regOut[8][2] ,
		\regOut[8][1] ,
		\regOut[8][0]  }),
	.FE_OFN4_write(FE_OFN21_write),
	.FE_OFN6_write(FE_OFN44_write),
	.FE_OFN34_write(FE_OFN34_write),
	.FE_OFN43_write(FE_OFN43_write),
	.clk__L2_N12(clk__L2_N12),
	.clk__L2_N2(clk__L2_N2),
	.clk__L2_N3(clk__L2_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   SingleReg_22 RegX_9 (
	.data({ \regIn[9][15] ,
		\regIn[9][14] ,
		\regIn[9][13] ,
		\regIn[9][12] ,
		\regIn[9][11] ,
		\regIn[9][10] ,
		\regIn[9][9] ,
		\regIn[9][8] ,
		\regIn[9][7] ,
		\regIn[9][6] ,
		\regIn[9][5] ,
		\regIn[9][4] ,
		\regIn[9][3] ,
		\regIn[9][2] ,
		\regIn[9][1] ,
		\regIn[9][0]  }),
	.clk(clk__L2_N0),
	.reset(reset),
	.write(FE_OFN21_write),
	.dataOut({ \regOut[9][15] ,
		\regOut[9][14] ,
		\regOut[9][13] ,
		\regOut[9][12] ,
		\regOut[9][11] ,
		\regOut[9][10] ,
		\regOut[9][9] ,
		\regOut[9][8] ,
		\regOut[9][7] ,
		\regOut[9][6] ,
		\regOut[9][5] ,
		\regOut[9][4] ,
		\regOut[9][3] ,
		\regOut[9][2] ,
		\regOut[9][1] ,
		\regOut[9][0]  }),
	.FE_OFN5_write(FE_OFN49_write),
	.FE_OFN6_write(FE_OFN44_write),
	.FE_OFN34_write(FE_OFN34_write),
	.FE_OFN47_write(FE_OFN47_write),
	.clk__L2_N12(clk__L2_N12),
	.clk__L2_N2(clk__L2_N2),
	.clk__L2_N3(clk__L2_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   SingleReg_21 RegX_10 (
	.data({ \regIn[10][15] ,
		\regIn[10][14] ,
		\regIn[10][13] ,
		\regIn[10][12] ,
		\regIn[10][11] ,
		\regIn[10][10] ,
		\regIn[10][9] ,
		\regIn[10][8] ,
		\regIn[10][7] ,
		\regIn[10][6] ,
		\regIn[10][5] ,
		\regIn[10][4] ,
		\regIn[10][3] ,
		\regIn[10][2] ,
		\regIn[10][1] ,
		\regIn[10][0]  }),
	.clk(clk__L2_N11),
	.reset(reset),
	.write(FE_OFN21_write),
	.dataOut({ \regOut[10][15] ,
		\regOut[10][14] ,
		\regOut[10][13] ,
		\regOut[10][12] ,
		\regOut[10][11] ,
		\regOut[10][10] ,
		\regOut[10][9] ,
		\regOut[10][8] ,
		\regOut[10][7] ,
		\regOut[10][6] ,
		\regOut[10][5] ,
		\regOut[10][4] ,
		\regOut[10][3] ,
		\regOut[10][2] ,
		\regOut[10][1] ,
		\regOut[10][0]  }),
	.FE_OFN6_write(FE_OFN44_write),
	.FE_OFN7_write(FE_OFN38_write),
	.FE_OFN9_write(FE_OFN55_write),
	.FE_OFN40_write(FE_OFN40_write),
	.FE_OFN43_write(FE_OFN43_write),
	.FE_OFN45_write(FE_OFN45_write),
	.FE_OFN50_write(FE_OFN50_write),
	.clk__L2_N12(clk__L2_N12), 
	.VDD(VDD), 
	.VSS(VSS));
   SingleReg_20 RegX_11 (
	.data({ \regIn[11][15] ,
		\regIn[11][14] ,
		\regIn[11][13] ,
		\regIn[11][12] ,
		\regIn[11][11] ,
		\regIn[11][10] ,
		\regIn[11][9] ,
		\regIn[11][8] ,
		\regIn[11][7] ,
		\regIn[11][6] ,
		\regIn[11][5] ,
		\regIn[11][4] ,
		\regIn[11][3] ,
		\regIn[11][2] ,
		\regIn[11][1] ,
		\regIn[11][0]  }),
	.clk(clk__L2_N11),
	.reset(reset),
	.write(FE_OFN21_write),
	.dataOut({ \regOut[11][15] ,
		\regOut[11][14] ,
		\regOut[11][13] ,
		\regOut[11][12] ,
		\regOut[11][11] ,
		\regOut[11][10] ,
		\regOut[11][9] ,
		\regOut[11][8] ,
		\regOut[11][7] ,
		\regOut[11][6] ,
		\regOut[11][5] ,
		\regOut[11][4] ,
		\regOut[11][3] ,
		\regOut[11][2] ,
		\regOut[11][1] ,
		\regOut[11][0]  }),
	.FE_OFN6_write(FE_OFN44_write),
	.FE_OFN7_write(FE_OFN38_write),
	.FE_OFN34_write(FE_OFN34_write),
	.FE_OFN38_write(FE_OFN38_write),
	.FE_OFN40_write(FE_OFN40_write),
	.FE_OFN43_write(FE_OFN43_write),
	.FE_OFN45_write(FE_OFN45_write),
	.clk__L2_N12(clk__L2_N12),
	.clk__L2_N2(clk__L2_N2),
	.clk__L2_N6(clk__L2_N6), 
	.VDD(VDD), 
	.VSS(VSS));
   SingleReg_19 RegX_12 (
	.data({ \regIn[12][15] ,
		\regIn[12][14] ,
		\regIn[12][13] ,
		\regIn[12][12] ,
		\regIn[12][11] ,
		\regIn[12][10] ,
		\regIn[12][9] ,
		\regIn[12][8] ,
		\regIn[12][7] ,
		\regIn[12][6] ,
		\regIn[12][5] ,
		\regIn[12][4] ,
		\regIn[12][3] ,
		\regIn[12][2] ,
		\regIn[12][1] ,
		\regIn[12][0]  }),
	.clk(clk__L2_N1),
	.reset(reset),
	.write(FE_OFN44_write),
	.dataOut({ \regOut[12][15] ,
		\regOut[12][14] ,
		\regOut[12][13] ,
		\regOut[12][12] ,
		\regOut[12][11] ,
		\regOut[12][10] ,
		\regOut[12][9] ,
		\regOut[12][8] ,
		\regOut[12][7] ,
		\regOut[12][6] ,
		\regOut[12][5] ,
		\regOut[12][4] ,
		\regOut[12][3] ,
		\regOut[12][2] ,
		\regOut[12][1] ,
		\regOut[12][0]  }),
	.FE_OFN7_write(FE_OFN38_write),
	.FE_OFN9_write(FE_OFN38_write),
	.FE_OFN50_write(FE_OFN50_write),
	.FE_OFN55_write(FE_OFN55_write),
	.clk__L2_N11(clk__L2_N11),
	.clk__L2_N12(clk__L2_N12),
	.clk__L2_N6(clk__L2_N6), 
	.VDD(VDD), 
	.VSS(VSS));
   SingleReg_18 RegX_13 (
	.data({ \regIn[13][15] ,
		\regIn[13][14] ,
		\regIn[13][13] ,
		\regIn[13][12] ,
		\regIn[13][11] ,
		\regIn[13][10] ,
		\regIn[13][9] ,
		\regIn[13][8] ,
		\regIn[13][7] ,
		\regIn[13][6] ,
		\regIn[13][5] ,
		\regIn[13][4] ,
		\regIn[13][3] ,
		\regIn[13][2] ,
		\regIn[13][1] ,
		\regIn[13][0]  }),
	.clk(clk__L2_N1),
	.reset(reset),
	.write(FE_OFN44_write),
	.dataOut({ \regOut[13][15] ,
		\regOut[13][14] ,
		\regOut[13][13] ,
		\regOut[13][12] ,
		\regOut[13][11] ,
		\regOut[13][10] ,
		\regOut[13][9] ,
		\regOut[13][8] ,
		\regOut[13][7] ,
		\regOut[13][6] ,
		\regOut[13][5] ,
		\regOut[13][4] ,
		\regOut[13][3] ,
		\regOut[13][2] ,
		\regOut[13][1] ,
		\regOut[13][0]  }),
	.FE_OFN7_write(FE_OFN38_write),
	.FE_OFN9_write(FE_OFN55_write),
	.FE_OFN50_write(FE_OFN50_write),
	.clk__L2_N11(clk__L2_N11),
	.clk__L2_N12(clk__L2_N12), 
	.VDD(VDD), 
	.VSS(VSS));
   SingleReg_17 RegX_14 (
	.data({ \regIn[14][15] ,
		\regIn[14][14] ,
		\regIn[14][13] ,
		\regIn[14][12] ,
		\regIn[14][11] ,
		\regIn[14][10] ,
		\regIn[14][9] ,
		\regIn[14][8] ,
		\regIn[14][7] ,
		\regIn[14][6] ,
		\regIn[14][5] ,
		\regIn[14][4] ,
		\regIn[14][3] ,
		\regIn[14][2] ,
		\regIn[14][1] ,
		\regIn[14][0]  }),
	.clk(clk__L2_N1),
	.reset(reset),
	.write(FE_OFN38_write),
	.dataOut({ \regOut[14][15] ,
		\regOut[14][14] ,
		\regOut[14][13] ,
		\regOut[14][12] ,
		\regOut[14][11] ,
		\regOut[14][10] ,
		\regOut[14][9] ,
		\regOut[14][8] ,
		\regOut[14][7] ,
		\regOut[14][6] ,
		\regOut[14][5] ,
		\regOut[14][4] ,
		\regOut[14][3] ,
		\regOut[14][2] ,
		\regOut[14][1] ,
		\regOut[14][0]  }),
	.FE_OFN9_write(FE_OFN55_write),
	.clk__L2_N11(clk__L2_N11), 
	.VDD(VDD), 
	.VSS(VSS));
   SingleReg_16 RegX_15 (
	.data({ \regIn[15][15] ,
		\regIn[15][14] ,
		\regIn[15][13] ,
		\regIn[15][12] ,
		\regIn[15][11] ,
		\regIn[15][10] ,
		\regIn[15][9] ,
		\regIn[15][8] ,
		\regIn[15][7] ,
		\regIn[15][6] ,
		\regIn[15][5] ,
		\regIn[15][4] ,
		\regIn[15][3] ,
		\regIn[15][2] ,
		\regIn[15][1] ,
		\regIn[15][0]  }),
	.clk(clk__L2_N1),
	.reset(reset),
	.write(FE_OFN44_write),
	.dataOut({ \regOut[15][15] ,
		\regOut[15][14] ,
		\regOut[15][13] ,
		\regOut[15][12] ,
		\regOut[15][11] ,
		\regOut[15][10] ,
		\regOut[15][9] ,
		\regOut[15][8] ,
		\regOut[15][7] ,
		\regOut[15][6] ,
		\regOut[15][5] ,
		\regOut[15][4] ,
		\regOut[15][3] ,
		\regOut[15][2] ,
		\regOut[15][1] ,
		\regOut[15][0]  }),
	.FE_OFN7_write(FE_OFN38_write),
	.FE_OFN9_write(FE_OFN55_write),
	.clk__L2_N11(clk__L2_N11), 
	.VDD(VDD), 
	.VSS(VSS));
   SingleReg_15 RegX_16 (
	.data({ \regIn[16][15] ,
		\regIn[16][14] ,
		\regIn[16][13] ,
		\regIn[16][12] ,
		\regIn[16][11] ,
		\regIn[16][10] ,
		\regIn[16][9] ,
		\regIn[16][8] ,
		\regIn[16][7] ,
		\regIn[16][6] ,
		\regIn[16][5] ,
		\regIn[16][4] ,
		\regIn[16][3] ,
		\regIn[16][2] ,
		\regIn[16][1] ,
		\regIn[16][0]  }),
	.clk(clk__L2_N10),
	.reset(reset),
	.write(FE_OFN18_write),
	.dataOut({ \regOut[16][15] ,
		\regOut[16][14] ,
		\regOut[16][13] ,
		\regOut[16][12] ,
		\regOut[16][11] ,
		\regOut[16][10] ,
		\regOut[16][9] ,
		\regOut[16][8] ,
		\regOut[16][7] ,
		\regOut[16][6] ,
		\regOut[16][5] ,
		\regOut[16][4] ,
		\regOut[16][3] ,
		\regOut[16][2] ,
		\regOut[16][1] ,
		\regOut[16][0]  }),
	.FE_OFN12_write(FE_OFN46_write),
	.FE_OFN3_write(FE_OFN18_write),
	.FE_OFN8_write(FE_OFN26_write),
	.FE_OFN26_write(FE_OFN26_write),
	.FE_OFN30_write(FE_OFN30_write),
	.clk__L2_N13(clk__L2_N13),
	.clk__L2_N4(clk__L2_N4),
	.clk__L2_N8(clk__L2_N8), 
	.VDD(VDD), 
	.VSS(VSS));
   SingleReg_14 RegX_17 (
	.data({ \regIn[17][15] ,
		\regIn[17][14] ,
		\regIn[17][13] ,
		\regIn[17][12] ,
		\regIn[17][11] ,
		\regIn[17][10] ,
		\regIn[17][9] ,
		\regIn[17][8] ,
		\regIn[17][7] ,
		\regIn[17][6] ,
		\regIn[17][5] ,
		\regIn[17][4] ,
		\regIn[17][3] ,
		\regIn[17][2] ,
		\regIn[17][1] ,
		\regIn[17][0]  }),
	.clk(clk__L2_N13),
	.reset(reset),
	.write(FE_OFN18_write),
	.dataOut({ \regOut[17][15] ,
		\regOut[17][14] ,
		\regOut[17][13] ,
		\regOut[17][12] ,
		\regOut[17][11] ,
		\regOut[17][10] ,
		\regOut[17][9] ,
		\regOut[17][8] ,
		\regOut[17][7] ,
		\regOut[17][6] ,
		\regOut[17][5] ,
		\regOut[17][4] ,
		\regOut[17][3] ,
		\regOut[17][2] ,
		\regOut[17][1] ,
		\regOut[17][0]  }),
	.FE_OFN10_write(FE_OFN46_write),
	.FE_OFN12_write(FE_OFN46_write),
	.FE_OFN3_write(FE_OFN26_write),
	.FE_OFN8_write(FE_OFN26_write),
	.FE_OFN30_write(FE_OFN30_write),
	.clk__L2_N4(clk__L2_N4),
	.clk__L2_N8(clk__L2_N8), 
	.VDD(VDD), 
	.VSS(VSS));
   SingleReg_13 RegX_18 (
	.data({ \regIn[18][15] ,
		\regIn[18][14] ,
		\regIn[18][13] ,
		\regIn[18][12] ,
		\regIn[18][11] ,
		\regIn[18][10] ,
		\regIn[18][9] ,
		\regIn[18][8] ,
		\regIn[18][7] ,
		\regIn[18][6] ,
		\regIn[18][5] ,
		\regIn[18][4] ,
		\regIn[18][3] ,
		\regIn[18][2] ,
		\regIn[18][1] ,
		\regIn[18][0]  }),
	.clk(clk__L2_N13),
	.reset(reset),
	.write(FE_OFN23_write),
	.dataOut({ \regOut[18][15] ,
		\regOut[18][14] ,
		\regOut[18][13] ,
		\regOut[18][12] ,
		\regOut[18][11] ,
		\regOut[18][10] ,
		\regOut[18][9] ,
		\regOut[18][8] ,
		\regOut[18][7] ,
		\regOut[18][6] ,
		\regOut[18][5] ,
		\regOut[18][4] ,
		\regOut[18][3] ,
		\regOut[18][2] ,
		\regOut[18][1] ,
		\regOut[18][0]  }),
	.FE_OFN3_write(FE_OFN18_write),
	.FE_OFN28_write(FE_OFN28_write),
	.clk__L2_N8(clk__L2_N8), 
	.VDD(VDD), 
	.VSS(VSS));
   SingleReg_12 RegX_19 (
	.data({ \regIn[19][15] ,
		\regIn[19][14] ,
		\regIn[19][13] ,
		\regIn[19][12] ,
		\regIn[19][11] ,
		\regIn[19][10] ,
		\regIn[19][9] ,
		\regIn[19][8] ,
		\regIn[19][7] ,
		\regIn[19][6] ,
		\regIn[19][5] ,
		\regIn[19][4] ,
		\regIn[19][3] ,
		\regIn[19][2] ,
		\regIn[19][1] ,
		\regIn[19][0]  }),
	.clk(clk__L2_N13),
	.reset(reset),
	.write(FE_OFN18_write),
	.dataOut({ \regOut[19][15] ,
		\regOut[19][14] ,
		\regOut[19][13] ,
		\regOut[19][12] ,
		\regOut[19][11] ,
		\regOut[19][10] ,
		\regOut[19][9] ,
		\regOut[19][8] ,
		\regOut[19][7] ,
		\regOut[19][6] ,
		\regOut[19][5] ,
		\regOut[19][4] ,
		\regOut[19][3] ,
		\regOut[19][2] ,
		\regOut[19][1] ,
		\regOut[19][0]  }),
	.FE_OFN12_write(FE_OFN46_write),
	.FE_OFN3_write(FE_OFN18_write),
	.FE_OFN23_write(FE_OFN23_write),
	.FE_OFN26_write(FE_OFN26_write),
	.FE_OFN28_write(FE_OFN28_write),
	.clk__L2_N8(clk__L2_N8), 
	.VDD(VDD), 
	.VSS(VSS));
   SingleReg_11 RegX_20 (
	.data({ \regIn[20][15] ,
		\regIn[20][14] ,
		\regIn[20][13] ,
		\regIn[20][12] ,
		\regIn[20][11] ,
		\regIn[20][10] ,
		\regIn[20][9] ,
		\regIn[20][8] ,
		\regIn[20][7] ,
		\regIn[20][6] ,
		\regIn[20][5] ,
		\regIn[20][4] ,
		\regIn[20][3] ,
		\regIn[20][2] ,
		\regIn[20][1] ,
		\regIn[20][0]  }),
	.clk(clk__L2_N0),
	.reset(reset),
	.write(FE_OFN48_write),
	.dataOut({ \regOut[20][15] ,
		\regOut[20][14] ,
		\regOut[20][13] ,
		\regOut[20][12] ,
		\regOut[20][11] ,
		\regOut[20][10] ,
		\regOut[20][9] ,
		\regOut[20][8] ,
		\regOut[20][7] ,
		\regOut[20][6] ,
		\regOut[20][5] ,
		\regOut[20][4] ,
		\regOut[20][3] ,
		\regOut[20][2] ,
		\regOut[20][1] ,
		\regOut[20][0]  }),
	.FE_OFN11_write(FE_OFN40_write),
	.FE_OFN5_write(FE_OFN40_write),
	.FE_OFN8_write(FE_OFN42_write),
	.FE_OFN49_write(FE_OFN49_write),
	.FE_OFN51_write(FE_OFN51_write),
	.FE_OFN53_write(FE_OFN53_write),
	.FE_OFN54_write(FE_OFN54_write),
	.FE_OFN56_write(FE_OFN56_write),
	.clk__L2_N10(clk__L2_N10),
	.clk__L2_N5(clk__L2_N5),
	.clk__L2_N6(clk__L2_N6), 
	.VDD(VDD), 
	.VSS(VSS));
   SingleReg_10 RegX_21 (
	.data({ \regIn[21][15] ,
		\regIn[21][14] ,
		\regIn[21][13] ,
		\regIn[21][12] ,
		\regIn[21][11] ,
		\regIn[21][10] ,
		\regIn[21][9] ,
		\regIn[21][8] ,
		\regIn[21][7] ,
		\regIn[21][6] ,
		\regIn[21][5] ,
		\regIn[21][4] ,
		\regIn[21][3] ,
		\regIn[21][2] ,
		\regIn[21][1] ,
		\regIn[21][0]  }),
	.clk(clk__L2_N0),
	.reset(reset),
	.write(FE_OFN26_write),
	.dataOut({ \regOut[21][15] ,
		\regOut[21][14] ,
		\regOut[21][13] ,
		\regOut[21][12] ,
		\regOut[21][11] ,
		\regOut[21][10] ,
		\regOut[21][9] ,
		\regOut[21][8] ,
		\regOut[21][7] ,
		\regOut[21][6] ,
		\regOut[21][5] ,
		\regOut[21][4] ,
		\regOut[21][3] ,
		\regOut[21][2] ,
		\regOut[21][1] ,
		\regOut[21][0]  }),
	.FE_OFN11_write(FE_OFN40_write),
	.FE_OFN4_write(FE_OFN47_write),
	.FE_OFN5_write(FE_OFN40_write),
	.FE_OFN8_write(FE_OFN42_write),
	.FE_OFN48_write(FE_OFN48_write),
	.FE_OFN49_write(FE_OFN49_write),
	.FE_OFN54_write(FE_OFN54_write),
	.FE_OFN56_write(FE_OFN56_write),
	.clk__L2_N10(clk__L2_N10),
	.clk__L2_N5(clk__L2_N5), 
	.VDD(VDD), 
	.VSS(VSS));
   SingleReg_9 RegX_22 (
	.data({ \regIn[22][15] ,
		\regIn[22][14] ,
		\regIn[22][13] ,
		\regIn[22][12] ,
		\regIn[22][11] ,
		\regIn[22][10] ,
		\regIn[22][9] ,
		\regIn[22][8] ,
		\regIn[22][7] ,
		\regIn[22][6] ,
		\regIn[22][5] ,
		\regIn[22][4] ,
		\regIn[22][3] ,
		\regIn[22][2] ,
		\regIn[22][1] ,
		\regIn[22][0]  }),
	.clk(clk__L2_N5),
	.reset(reset),
	.write(FE_OFN40_write),
	.dataOut({ \regOut[22][15] ,
		\regOut[22][14] ,
		\regOut[22][13] ,
		\regOut[22][12] ,
		\regOut[22][11] ,
		\regOut[22][10] ,
		\regOut[22][9] ,
		\regOut[22][8] ,
		\regOut[22][7] ,
		\regOut[22][6] ,
		\regOut[22][5] ,
		\regOut[22][4] ,
		\regOut[22][3] ,
		\regOut[22][2] ,
		\regOut[22][1] ,
		\regOut[22][0]  }),
	.FE_OFN13_write(FE_OFN40_write),
	.FE_OFN5_write(FE_OFN51_write),
	.FE_OFN56_write(FE_OFN56_write),
	.FE_OFN57_write(FE_OFN57_write),
	.FE_OFN58_write(FE_OFN58_write),
	.clk__L2_N6(clk__L2_N6),
	.clk__L2_N9(clk__L2_N9), 
	.VDD(VDD), 
	.VSS(VSS));
   SingleReg_8 RegX_23 (
	.data({ \regIn[23][15] ,
		\regIn[23][14] ,
		\regIn[23][13] ,
		\regIn[23][12] ,
		\regIn[23][11] ,
		\regIn[23][10] ,
		\regIn[23][9] ,
		\regIn[23][8] ,
		\regIn[23][7] ,
		\regIn[23][6] ,
		\regIn[23][5] ,
		\regIn[23][4] ,
		\regIn[23][3] ,
		\regIn[23][2] ,
		\regIn[23][1] ,
		\regIn[23][0]  }),
	.clk(clk__L2_N0),
	.reset(reset),
	.write(FE_OFN40_write),
	.dataOut({ \regOut[23][15] ,
		\regOut[23][14] ,
		\regOut[23][13] ,
		\regOut[23][12] ,
		\regOut[23][11] ,
		\regOut[23][10] ,
		\regOut[23][9] ,
		\regOut[23][8] ,
		\regOut[23][7] ,
		\regOut[23][6] ,
		\regOut[23][5] ,
		\regOut[23][4] ,
		\regOut[23][3] ,
		\regOut[23][2] ,
		\regOut[23][1] ,
		\regOut[23][0]  }),
	.FE_OFN13_write(FE_OFN57_write),
	.FE_OFN5_write(FE_OFN40_write),
	.FE_OFN8_write(FE_OFN42_write),
	.FE_OFN53_write(FE_OFN53_write),
	.FE_OFN54_write(FE_OFN54_write),
	.FE_OFN56_write(FE_OFN56_write),
	.clk__L2_N5(clk__L2_N5),
	.clk__L2_N6(clk__L2_N6), 
	.VDD(VDD), 
	.VSS(VSS));
   SingleReg_7 RegX_24 (
	.data({ \regIn[24][15] ,
		\regIn[24][14] ,
		\regIn[24][13] ,
		\regIn[24][12] ,
		\regIn[24][11] ,
		\regIn[24][10] ,
		\regIn[24][9] ,
		\regIn[24][8] ,
		\regIn[24][7] ,
		\regIn[24][6] ,
		\regIn[24][5] ,
		\regIn[24][4] ,
		\regIn[24][3] ,
		\regIn[24][2] ,
		\regIn[24][1] ,
		\regIn[24][0]  }),
	.clk(clk__L2_N0),
	.reset(reset),
	.write(FE_OFN26_write),
	.dataOut({ \regOut[24][15] ,
		\regOut[24][14] ,
		\regOut[24][13] ,
		\regOut[24][12] ,
		\regOut[24][11] ,
		\regOut[24][10] ,
		\regOut[24][9] ,
		\regOut[24][8] ,
		\regOut[24][7] ,
		\regOut[24][6] ,
		\regOut[24][5] ,
		\regOut[24][4] ,
		\regOut[24][3] ,
		\regOut[24][2] ,
		\regOut[24][1] ,
		\regOut[24][0]  }),
	.FE_OFN11_write(FE_OFN54_write),
	.FE_OFN5_write(FE_OFN49_write),
	.FE_OFN8_write(FE_OFN26_write),
	.FE_OFN42_write(FE_OFN42_write),
	.FE_OFN46_write(FE_OFN46_write),
	.FE_OFN48_write(FE_OFN48_write),
	.clk__L2_N10(clk__L2_N10),
	.clk__L2_N4(clk__L2_N4), 
	.VDD(VDD), 
	.VSS(VSS));
   SingleReg_6 RegX_25 (
	.data({ \regIn[25][15] ,
		\regIn[25][14] ,
		\regIn[25][13] ,
		\regIn[25][12] ,
		\regIn[25][11] ,
		\regIn[25][10] ,
		\regIn[25][9] ,
		\regIn[25][8] ,
		\regIn[25][7] ,
		\regIn[25][6] ,
		\regIn[25][5] ,
		\regIn[25][4] ,
		\regIn[25][3] ,
		\regIn[25][2] ,
		\regIn[25][1] ,
		\regIn[25][0]  }),
	.clk(clk__L2_N0),
	.reset(reset),
	.write(FE_OFN26_write),
	.dataOut({ \regOut[25][15] ,
		\regOut[25][14] ,
		\regOut[25][13] ,
		\regOut[25][12] ,
		\regOut[25][11] ,
		\regOut[25][10] ,
		\regOut[25][9] ,
		\regOut[25][8] ,
		\regOut[25][7] ,
		\regOut[25][6] ,
		\regOut[25][5] ,
		\regOut[25][4] ,
		\regOut[25][3] ,
		\regOut[25][2] ,
		\regOut[25][1] ,
		\regOut[25][0]  }),
	.FE_OFN5_write(FE_OFN49_write),
	.FE_OFN8_write(FE_OFN26_write),
	.FE_OFN42_write(FE_OFN42_write),
	.FE_OFN46_write(FE_OFN46_write),
	.FE_OFN48_write(FE_OFN48_write),
	.clk__L2_N10(clk__L2_N10),
	.clk__L2_N4(clk__L2_N4), 
	.VDD(VDD), 
	.VSS(VSS));
   SingleReg_5 RegX_26 (
	.data({ \regIn[26][15] ,
		\regIn[26][14] ,
		\regIn[26][13] ,
		\regIn[26][12] ,
		\regIn[26][11] ,
		\regIn[26][10] ,
		\regIn[26][9] ,
		\regIn[26][8] ,
		\regIn[26][7] ,
		\regIn[26][6] ,
		\regIn[26][5] ,
		\regIn[26][4] ,
		\regIn[26][3] ,
		\regIn[26][2] ,
		\regIn[26][1] ,
		\regIn[26][0]  }),
	.clk(clk__L2_N10),
	.reset(reset),
	.write(FE_OFN46_write),
	.dataOut({ \regOut[26][15] ,
		\regOut[26][14] ,
		\regOut[26][13] ,
		\regOut[26][12] ,
		\regOut[26][11] ,
		\regOut[26][10] ,
		\regOut[26][9] ,
		\regOut[26][8] ,
		\regOut[26][7] ,
		\regOut[26][6] ,
		\regOut[26][5] ,
		\regOut[26][4] ,
		\regOut[26][3] ,
		\regOut[26][2] ,
		\regOut[26][1] ,
		\regOut[26][0]  }),
	.FE_OFN1_write(FE_OFN25_write),
	.FE_OFN8_write(FE_OFN26_write),
	.FE_OFN35_write(FE_OFN35_write),
	.FE_OFN39_write(FE_OFN39_write),
	.clk__L2_N4(clk__L2_N4), 
	.VDD(VDD), 
	.VSS(VSS));
   SingleReg_4 RegX_27 (
	.data({ \regIn[27][15] ,
		\regIn[27][14] ,
		\regIn[27][13] ,
		\regIn[27][12] ,
		\regIn[27][11] ,
		\regIn[27][10] ,
		\regIn[27][9] ,
		\regIn[27][8] ,
		\regIn[27][7] ,
		\regIn[27][6] ,
		\regIn[27][5] ,
		\regIn[27][4] ,
		\regIn[27][3] ,
		\regIn[27][2] ,
		\regIn[27][1] ,
		\regIn[27][0]  }),
	.clk(clk__L2_N10),
	.reset(reset),
	.write(FE_OFN46_write),
	.dataOut({ \regOut[27][15] ,
		\regOut[27][14] ,
		\regOut[27][13] ,
		\regOut[27][12] ,
		\regOut[27][11] ,
		\regOut[27][10] ,
		\regOut[27][9] ,
		\regOut[27][8] ,
		\regOut[27][7] ,
		\regOut[27][6] ,
		\regOut[27][5] ,
		\regOut[27][4] ,
		\regOut[27][3] ,
		\regOut[27][2] ,
		\regOut[27][1] ,
		\regOut[27][0]  }),
	.FE_OFN8_write(FE_OFN26_write),
	.FE_OFN35_write(FE_OFN35_write),
	.FE_OFN39_write(FE_OFN39_write),
	.clk__L2_N13(clk__L2_N13),
	.clk__L2_N4(clk__L2_N4), 
	.VDD(VDD), 
	.VSS(VSS));
   SingleReg_3 RegX_28 (
	.data({ \regIn[28][15] ,
		\regIn[28][14] ,
		\regIn[28][13] ,
		\regIn[28][12] ,
		\regIn[28][11] ,
		\regIn[28][10] ,
		\regIn[28][9] ,
		\regIn[28][8] ,
		\regIn[28][7] ,
		\regIn[28][6] ,
		\regIn[28][5] ,
		\regIn[28][4] ,
		\regIn[28][3] ,
		\regIn[28][2] ,
		\regIn[28][1] ,
		\regIn[28][0]  }),
	.clk(clk__L2_N1),
	.reset(reset),
	.write(FE_OFN59_write),
	.dataOut({ \regOut[28][15] ,
		\regOut[28][14] ,
		\regOut[28][13] ,
		\regOut[28][12] ,
		\regOut[28][11] ,
		\regOut[28][10] ,
		\regOut[28][9] ,
		\regOut[28][8] ,
		\regOut[28][7] ,
		\regOut[28][6] ,
		\regOut[28][5] ,
		\regOut[28][4] ,
		\regOut[28][3] ,
		\regOut[28][2] ,
		\regOut[28][1] ,
		\regOut[28][0]  }),
	.FE_OFN14_write(FE_OFN58_write),
	.FE_OFN9_write(FE_OFN55_write),
	.clk__L2_N6(clk__L2_N6),
	.clk__L2_N9(clk__L2_N9), 
	.VDD(VDD), 
	.VSS(VSS));
   SingleReg_2 RegX_29 (
	.data({ \regIn[29][15] ,
		\regIn[29][14] ,
		\regIn[29][13] ,
		\regIn[29][12] ,
		\regIn[29][11] ,
		\regIn[29][10] ,
		\regIn[29][9] ,
		\regIn[29][8] ,
		\regIn[29][7] ,
		\regIn[29][6] ,
		\regIn[29][5] ,
		\regIn[29][4] ,
		\regIn[29][3] ,
		\regIn[29][2] ,
		\regIn[29][1] ,
		\regIn[29][0]  }),
	.clk(clk__L2_N1),
	.reset(reset),
	.write(FE_OFN59_write),
	.dataOut({ \regOut[29][15] ,
		\regOut[29][14] ,
		\regOut[29][13] ,
		\regOut[29][12] ,
		\regOut[29][11] ,
		\regOut[29][10] ,
		\regOut[29][9] ,
		\regOut[29][8] ,
		\regOut[29][7] ,
		\regOut[29][6] ,
		\regOut[29][5] ,
		\regOut[29][4] ,
		\regOut[29][3] ,
		\regOut[29][2] ,
		\regOut[29][1] ,
		\regOut[29][0]  }),
	.FE_OFN14_write(FE_OFN58_write),
	.clk__L2_N6(clk__L2_N6),
	.clk__L2_N9(clk__L2_N9), 
	.VDD(VDD), 
	.VSS(VSS));
   SingleReg_1 RegX_30 (
	.data({ \regIn[30][15] ,
		\regIn[30][14] ,
		\regIn[30][13] ,
		\regIn[30][12] ,
		\regIn[30][11] ,
		\regIn[30][10] ,
		\regIn[30][9] ,
		\regIn[30][8] ,
		\regIn[30][7] ,
		\regIn[30][6] ,
		\regIn[30][5] ,
		\regIn[30][4] ,
		\regIn[30][3] ,
		\regIn[30][2] ,
		\regIn[30][1] ,
		\regIn[30][0]  }),
	.clk(clk__L2_N6),
	.reset(reset),
	.write(FE_OFN56_write),
	.dataOut({ \regOut[30][15] ,
		\regOut[30][14] ,
		\regOut[30][13] ,
		\regOut[30][12] ,
		\regOut[30][11] ,
		\regOut[30][10] ,
		\regOut[30][9] ,
		\regOut[30][8] ,
		\regOut[30][7] ,
		\regOut[30][6] ,
		\regOut[30][5] ,
		\regOut[30][4] ,
		\regOut[30][3] ,
		\regOut[30][2] ,
		\regOut[30][1] ,
		\regOut[30][0]  }),
	.FE_OFN13_write(FE_OFN40_write),
	.FE_OFN14_write(FE_OFN58_write),
	.FE_OFN57_write(FE_OFN57_write),
	.FE_OFN58_write(FE_OFN58_write),
	.FE_OFN59_write(FE_OFN59_write),
	.clk__L2_N9(clk__L2_N9), 
	.VDD(VDD), 
	.VSS(VSS));
   SingleReg_0 RegX_31 (
	.data({ \regIn[31][15] ,
		\regIn[31][14] ,
		\regIn[31][13] ,
		\regIn[31][12] ,
		\regIn[31][11] ,
		\regIn[31][10] ,
		\regIn[31][9] ,
		\regIn[31][8] ,
		\regIn[31][7] ,
		\regIn[31][6] ,
		\regIn[31][5] ,
		\regIn[31][4] ,
		\regIn[31][3] ,
		\regIn[31][2] ,
		\regIn[31][1] ,
		\regIn[31][0]  }),
	.clk(clk__L2_N1),
	.reset(reset),
	.write(FE_OFN56_write),
	.dataOut({ \regOut[31][15] ,
		\regOut[31][14] ,
		\regOut[31][13] ,
		\regOut[31][12] ,
		\regOut[31][11] ,
		\regOut[31][10] ,
		\regOut[31][9] ,
		\regOut[31][8] ,
		\regOut[31][7] ,
		\regOut[31][6] ,
		\regOut[31][5] ,
		\regOut[31][4] ,
		\regOut[31][3] ,
		\regOut[31][2] ,
		\regOut[31][1] ,
		\regOut[31][0]  }),
	.FE_OFN13_write(FE_OFN40_write),
	.FE_OFN14_write(FE_OFN58_write),
	.FE_OFN9_write(FE_OFN55_write),
	.FE_OFN57_write(FE_OFN57_write),
	.FE_OFN58_write(FE_OFN58_write),
	.FE_OFN59_write(FE_OFN59_write),
	.clk__L2_N6(clk__L2_N6),
	.clk__L2_N9(clk__L2_N9), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUF_X1 U1789 (
	.Z(n1271),
	.A(N208), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2_X1 U1811 (
	.ZN(N326),
	.A2(N307),
	.A1(addressIn[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2_X1 U1812 (
	.ZN(N302),
	.A2(N307),
	.A1(addressIn[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2_X1 U1813 (
	.ZN(N320),
	.A2(N307),
	.A1(addressIn[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2_X1 U1814 (
	.ZN(N296),
	.A2(N307),
	.A1(addressIn[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2_X1 U1815 (
	.ZN(N338),
	.A2(N307),
	.A1(addressIn[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2_X1 U1816 (
	.ZN(N314),
	.A2(N307),
	.A1(addressIn[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2_X1 U1817 (
	.ZN(N332),
	.A2(N307),
	.A1(addressIn[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1818 (
	.ZN(N245),
	.A(addressIn[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2_X1 U1819 (
	.ZN(N308),
	.A2(N307),
	.A1(addressIn[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2_X1 U1822 (
	.ZN(N254),
	.A2(N253),
	.A1(addressIn[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2_X1 U1823 (
	.ZN(N351),
	.A2(N386),
	.A1(addressIn[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2_X1 U1824 (
	.ZN(N303),
	.A2(N302),
	.A1(addressIn[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2_X1 U1825 (
	.ZN(N203),
	.A2(N202),
	.A1(addressIn[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2_X1 U1826 (
	.ZN(N196),
	.A2(N195),
	.A1(addressIn[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2_X1 U1827 (
	.ZN(N248),
	.A2(N247),
	.A1(addressIn[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2_X1 U1828 (
	.ZN(N297),
	.A2(N296),
	.A1(addressIn[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2_X1 U1829 (
	.ZN(N345),
	.A2(N386),
	.A1(addressIn[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2_X1 U1830 (
	.ZN(N363),
	.A2(N386),
	.A1(addressIn[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2_X1 U1831 (
	.ZN(N216),
	.A2(N215),
	.A1(addressIn[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2_X1 U1832 (
	.ZN(N315),
	.A2(N314),
	.A1(addressIn[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2_X1 U1833 (
	.ZN(N266),
	.A2(N265),
	.A1(addressIn[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2_X1 U1834 (
	.ZN(N357),
	.A2(N386),
	.A1(addressIn[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2_X1 U1835 (
	.ZN(N210),
	.A2(N209),
	.A1(addressIn[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2_X1 U1836 (
	.ZN(N260),
	.A2(N259),
	.A1(addressIn[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2_X1 U1837 (
	.ZN(N309),
	.A2(N308),
	.A1(addressIn[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1838 (
	.ZN(N220),
	.A(addressIn[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2_X1 U1841 (
	.ZN(N255),
	.A2(N254),
	.A1(addressIn[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2_X1 U1842 (
	.ZN(N352),
	.A2(N351),
	.A1(addressIn[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2_X1 U1843 (
	.ZN(N230),
	.A2(N229),
	.A1(addressIn[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2_X1 U1844 (
	.ZN(N304),
	.A2(N303),
	.A1(addressIn[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2_X1 U1845 (
	.ZN(N328),
	.A2(N327),
	.A1(addressIn[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2_X1 U1846 (
	.ZN(N204),
	.A2(N203),
	.A1(addressIn[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2_X1 U1847 (
	.ZN(N279),
	.A2(N278),
	.A1(addressIn[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2_X1 U1848 (
	.ZN(N197),
	.A2(N196),
	.A1(addressIn[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2_X1 U1849 (
	.ZN(N224),
	.A2(N223),
	.A1(addressIn[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2_X1 U1850 (
	.ZN(N273),
	.A2(N272),
	.A1(addressIn[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2_X1 U1851 (
	.ZN(N298),
	.A2(N297),
	.A1(addressIn[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2_X1 U1852 (
	.ZN(N322),
	.A2(N321),
	.A1(addressIn[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2_X1 U1853 (
	.ZN(N249),
	.A2(N248),
	.A1(addressIn[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2_X1 U1854 (
	.ZN(N346),
	.A2(N345),
	.A1(addressIn[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2_X1 U1855 (
	.ZN(N376),
	.A2(N387),
	.A1(addressIn[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2_X1 U1856 (
	.ZN(N370),
	.A2(N387),
	.A1(addressIn[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1857 (
	.ZN(N207),
	.A(addressIn[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2_X1 U1860 (
	.ZN(N198),
	.A2(N197),
	.A1(addressIn[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2_X1 U1861 (
	.ZN(N383),
	.A2(N388),
	.A1(addressIn[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2_X1 U1862 (
	.ZN(N250),
	.A2(N249),
	.A1(addressIn[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2_X1 U1863 (
	.ZN(N347),
	.A2(N346),
	.A1(addressIn[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2_X1 U1864 (
	.ZN(N274),
	.A2(N273),
	.A1(addressIn[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2_X1 U1865 (
	.ZN(N225),
	.A2(N224),
	.A1(addressIn[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2_X1 U1866 (
	.ZN(N299),
	.A2(N298),
	.A1(addressIn[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2_X1 U1867 (
	.ZN(N323),
	.A2(N322),
	.A1(addressIn[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2_X1 U1868 (
	.ZN(N359),
	.A2(N358),
	.A1(addressIn[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2_X1 U1869 (
	.ZN(N371),
	.A2(N370),
	.A1(addressIn[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2_X1 U1870 (
	.ZN(N335),
	.A2(N334),
	.A1(addressIn[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2_X1 U1871 (
	.ZN(N212),
	.A2(N211),
	.A1(addressIn[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2_X1 U1872 (
	.ZN(N311),
	.A2(N310),
	.A1(addressIn[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2_X1 U1873 (
	.ZN(N262),
	.A2(N261),
	.A1(addressIn[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2_X1 U1874 (
	.ZN(N237),
	.A2(N236),
	.A1(addressIn[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2_X1 U1875 (
	.ZN(N286),
	.A2(N285),
	.A1(addressIn[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   INV_X1 U1876 (
	.ZN(N200),
	.A(addressIn[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2_X1 U1878 (
	.ZN(N253),
	.A2(n1271),
	.A1(N245), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2_X1 U1879 (
	.ZN(N277),
	.A2(n1271),
	.A1(N245), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2_X1 U1880 (
	.ZN(N228),
	.A2(n1271),
	.A1(addressIn[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2_X1 U1881 (
	.ZN(N271),
	.A2(n1271),
	.A1(N245), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2_X1 U1882 (
	.ZN(N202),
	.A2(n1271),
	.A1(addressIn[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2_X1 U1883 (
	.ZN(N222),
	.A2(n1271),
	.A1(addressIn[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2_X1 U1884 (
	.ZN(N247),
	.A2(n1271),
	.A1(N245), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2_X1 U1885 (
	.ZN(N195),
	.A2(n1271),
	.A1(addressIn[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2_X1 U1886 (
	.ZN(N289),
	.A2(n1271),
	.A1(N245), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2_X1 U1887 (
	.ZN(N240),
	.A2(n1271),
	.A1(addressIn[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2_X1 U1888 (
	.ZN(N265),
	.A2(n1271),
	.A1(N245), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2_X1 U1889 (
	.ZN(N283),
	.A2(n1271),
	.A1(N245), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2_X1 U1890 (
	.ZN(N215),
	.A2(n1271),
	.A1(addressIn[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2_X1 U1891 (
	.ZN(N234),
	.A2(n1271),
	.A1(addressIn[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2_X1 U1892 (
	.ZN(N259),
	.A2(n1271),
	.A1(N245), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2_X1 U1893 (
	.ZN(N209),
	.A2(n1271),
	.A1(addressIn[3]), 
	.VDD(VDD), 
	.VSS(VSS));

   // Fillers and physical instances.
   FILLCELL_X2 FILL_1085 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_1084 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_1083 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X4 FILL_1082 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X8 FILL_1081 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X32 FILL_1080 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X8 FILL_1079 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_1078 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X4 FILL_1077 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_1076 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X8 FILL_1075 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_1074 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X4 FILL_1073 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_1072 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_1071 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_1070 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X4 FILL_1069 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X16 FILL_1068 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_1067 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_1066 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_1065 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_1064 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_1063 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X4 FILL_1062 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_1061 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_1060 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X4 FILL_1059 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_1058 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_1057 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_1056 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_1055 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_1054 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_1053 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_1052 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X32 FILL_1051 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X32 FILL_1050 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X4 FILL_1049 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_1048 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_1047 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_1046 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X4 FILL_1045 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_1044 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_1043 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X4 FILL_1042 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X8 FILL_1041 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_1040 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_1039 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X4 FILL_1038 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X8 FILL_1037 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_1036 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_1035 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_1034 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X4 FILL_1033 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_1032 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_1031 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_1030 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X4 FILL_1029 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X32 FILL_1028 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_1027 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_1026 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_1025 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_1024 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X4 FILL_1023 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X4 FILL_1022 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_1021 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_1020 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_1019 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_1018 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_1017 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_1016 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X4 FILL_1015 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_1014 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X4 FILL_1013 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X8 FILL_1012 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_1011 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_1010 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_1009 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X4 FILL_1008 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_1007 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_1006 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_1005 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_1004 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X32 FILL_1003 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_1002 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X8 FILL_1001 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X32 FILL_1000 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_999 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_998 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_997 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_996 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_995 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_994 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X4 FILL_993 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X4 FILL_992 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_991 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_990 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X4 FILL_989 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_988 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_987 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_986 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_985 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X4 FILL_984 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_983 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_982 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_981 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X4 FILL_980 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_979 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_978 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X8 FILL_977 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_976 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X8 FILL_975 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_974 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_973 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_972 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_971 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_970 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_969 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_968 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_967 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_966 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_965 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X4 FILL_964 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_963 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_962 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_961 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X4 FILL_960 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X16 FILL_959 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_958 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_957 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_956 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X8 FILL_955 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X16 FILL_954 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_953 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_952 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_951 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_950 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X4 FILL_949 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_948 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_947 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X4 FILL_946 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_945 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X4 FILL_944 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_943 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_942 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_941 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X4 FILL_940 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_939 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_938 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_937 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X4 FILL_936 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_935 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_934 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_933 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X4 FILL_932 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_931 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_930 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X4 FILL_929 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X4 FILL_928 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X8 FILL_927 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X32 FILL_926 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_925 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X4 FILL_924 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_923 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X8 FILL_922 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X32 FILL_921 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_920 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_919 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_918 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X4 FILL_917 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X16 FILL_916 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_915 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_914 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_913 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_912 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X4 FILL_911 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_910 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_909 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_908 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_907 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X8 FILL_906 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_905 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_904 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_903 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_902 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_901 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_900 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_899 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_898 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_897 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_896 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_895 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X8 FILL_894 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_893 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_892 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X32 FILL_891 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_890 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_889 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_888 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X8 FILL_887 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_886 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X4 FILL_885 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X4 FILL_884 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_883 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_882 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X8 FILL_881 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_880 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X8 FILL_879 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_878 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_877 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_876 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_875 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_874 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_873 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_872 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_871 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_870 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_869 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_868 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_867 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X16 FILL_866 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X32 FILL_865 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_864 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_863 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_862 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_861 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_860 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_859 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X4 FILL_858 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_857 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_856 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_855 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_854 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X4 FILL_853 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X16 FILL_852 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_851 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X8 FILL_850 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_849 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_848 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_847 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_846 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_845 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X8 FILL_844 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X8 FILL_843 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X16 FILL_842 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_841 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_840 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_839 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_838 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_837 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_836 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_835 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_834 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_833 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_832 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_831 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_830 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_829 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X4 FILL_828 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X16 FILL_827 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_826 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X4 FILL_825 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_824 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_823 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_822 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X4 FILL_821 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_820 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_819 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_818 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_817 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X32 FILL_816 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X4 FILL_815 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_814 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_813 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_812 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X4 FILL_811 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_810 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_809 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X8 FILL_808 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_807 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X4 FILL_806 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_805 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_804 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_803 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_802 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_801 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_800 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X4 FILL_799 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_798 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_797 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_796 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X4 FILL_795 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_794 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_793 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_792 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_791 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_790 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_789 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_788 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_787 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_786 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_785 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_784 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_783 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X4 FILL_782 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_781 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_780 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_779 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_778 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_777 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_776 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_775 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_774 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X8 FILL_773 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_772 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_771 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_770 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_769 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_768 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X4 FILL_767 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_766 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_765 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_764 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_763 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X8 FILL_762 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_761 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_760 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_759 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X4 FILL_758 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_757 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_756 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_755 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X4 FILL_754 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_753 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_752 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_751 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_750 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X4 FILL_749 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_748 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_747 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_746 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_745 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_744 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_743 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_742 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X4 FILL_741 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X4 FILL_740 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_739 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_738 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_737 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_736 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_735 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_734 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X8 FILL_733 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_732 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_731 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_730 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X8 FILL_729 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_728 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X4 FILL_727 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_726 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_725 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_724 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X4 FILL_723 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_722 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_721 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_720 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_719 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_718 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X4 FILL_717 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_716 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_715 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_714 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_713 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X8 FILL_712 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_711 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_710 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_709 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_708 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_707 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X4 FILL_706 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_705 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_704 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_703 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_702 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_701 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_700 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_699 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_698 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_697 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_696 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_695 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_694 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_693 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_692 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_691 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_690 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_689 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_688 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_687 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_686 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_685 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_684 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_683 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X4 FILL_682 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_681 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_680 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_679 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X4 FILL_678 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X4 FILL_677 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_676 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X8 FILL_675 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_674 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_673 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_672 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_671 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X4 FILL_670 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_669 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_668 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_667 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X4 FILL_666 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_665 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_664 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_663 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_662 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_661 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_660 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X4 FILL_659 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_658 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X4 FILL_657 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X8 FILL_656 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_655 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_654 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_653 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_652 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_651 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_650 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_649 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_648 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_647 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_646 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_645 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_644 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X4 FILL_643 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_642 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_641 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X4 FILL_640 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_639 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X4 FILL_638 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_637 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_636 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X4 FILL_635 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_634 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_633 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_632 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_631 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_630 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_629 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X4 FILL_628 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_627 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_626 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_625 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X4 FILL_624 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_623 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X4 FILL_622 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_621 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_620 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_619 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_618 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_617 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_616 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X4 FILL_615 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_614 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X8 FILL_613 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_612 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_611 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_610 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_609 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_608 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_607 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_606 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_605 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X16 FILL_604 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X4 FILL_603 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_602 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X4 FILL_601 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_600 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_599 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X4 FILL_598 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_597 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_596 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X4 FILL_595 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_594 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_593 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_592 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_591 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_590 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_589 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_588 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_587 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_586 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_585 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X4 FILL_584 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_583 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_582 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_581 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_580 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_579 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_578 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_577 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_576 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_575 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_574 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_573 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_572 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_571 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_570 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_569 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X4 FILL_568 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_567 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_566 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_565 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_564 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_563 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_562 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_561 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_560 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_559 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X8 FILL_558 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X8 FILL_557 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_556 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_555 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_554 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_553 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_552 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X4 FILL_551 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X8 FILL_550 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X32 FILL_549 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X4 FILL_548 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X4 FILL_547 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_546 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_545 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_544 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X4 FILL_543 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_542 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X4 FILL_541 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_540 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_539 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_538 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_537 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_536 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_535 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_534 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_533 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_532 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_531 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_530 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_529 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X4 FILL_528 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_527 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_526 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_525 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X4 FILL_524 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_523 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_522 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X4 FILL_521 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_520 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X4 FILL_519 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_518 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X4 FILL_517 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_516 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_515 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_514 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_513 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_512 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_511 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_510 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_509 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_508 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_507 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_506 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X4 FILL_505 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_504 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_503 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_502 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X8 FILL_501 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_500 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_499 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_498 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_497 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X4 FILL_496 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_495 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_494 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X4 FILL_493 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_492 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_491 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_490 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X4 FILL_489 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X8 FILL_488 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_487 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_486 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_485 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X4 FILL_484 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_483 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_482 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X4 FILL_481 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_480 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_479 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_478 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_477 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_476 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_475 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_474 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_473 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X4 FILL_472 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_471 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_470 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_469 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X4 FILL_468 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X16 FILL_467 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_466 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X4 FILL_465 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_464 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_463 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_462 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X4 FILL_461 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X8 FILL_460 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_459 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_458 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_457 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_456 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X4 FILL_455 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_454 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_453 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X4 FILL_452 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_451 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_450 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_449 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X4 FILL_448 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X8 FILL_447 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_446 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_445 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_444 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_443 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_442 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X4 FILL_441 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_440 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_439 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X8 FILL_438 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_437 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_436 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_435 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_434 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X4 FILL_433 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_432 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_431 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_430 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_429 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_428 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X4 FILL_427 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_426 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_425 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_424 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X4 FILL_423 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_422 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_421 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_420 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X4 FILL_419 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_418 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X4 FILL_417 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_416 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_415 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_414 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_413 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_412 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_411 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_410 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X4 FILL_409 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_408 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_407 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_406 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_405 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X8 FILL_404 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_403 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_402 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_401 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_400 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_399 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_398 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_397 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_396 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_395 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_394 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_393 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_392 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_391 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_390 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_389 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_388 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_387 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_386 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X4 FILL_385 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_384 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_383 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_382 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_381 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X4 FILL_380 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_379 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_378 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_377 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_376 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X4 FILL_375 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_374 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X4 FILL_373 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X8 FILL_372 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_371 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X4 FILL_370 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_369 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_368 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_367 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_366 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_365 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_364 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_363 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_362 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_361 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X4 FILL_360 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X4 FILL_359 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X8 FILL_358 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_357 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_356 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_355 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X4 FILL_354 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X8 FILL_353 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_352 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_351 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_350 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_349 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_348 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_347 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_346 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_345 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X4 FILL_344 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_343 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_342 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_341 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_340 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_339 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_338 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_337 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_336 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_335 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_334 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_333 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_332 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_331 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_330 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_329 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X4 FILL_328 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X16 FILL_327 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_326 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X4 FILL_325 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_324 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_323 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_322 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_321 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_320 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_319 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_318 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_317 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_316 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_315 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_314 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_313 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_312 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_311 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_310 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X4 FILL_309 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_308 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_307 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_306 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_305 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_304 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_303 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_302 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_301 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X4 FILL_300 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_299 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_298 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_297 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X8 FILL_296 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X4 FILL_295 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_294 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_293 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_292 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_291 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_290 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_289 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X8 FILL_288 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X4 FILL_287 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_286 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_285 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_284 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_283 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_282 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_281 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_280 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_279 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_278 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_277 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_276 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_275 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_274 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X4 FILL_273 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_272 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X4 FILL_271 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_270 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_269 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_268 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_267 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X16 FILL_266 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_265 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X4 FILL_264 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_263 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_262 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_261 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_260 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X8 FILL_259 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_258 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X4 FILL_257 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_256 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_255 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X8 FILL_254 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X4 FILL_253 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_252 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X4 FILL_251 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_250 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_249 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_248 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_247 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_246 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_245 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_244 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X4 FILL_243 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_242 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X4 FILL_241 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X4 FILL_240 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_239 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_238 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_237 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_236 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X8 FILL_235 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_234 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_233 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_232 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X4 FILL_231 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X8 FILL_230 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_229 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_228 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X8 FILL_227 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_226 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_225 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_224 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_223 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_222 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_221 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_220 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_219 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_218 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_217 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_216 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X4 FILL_215 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_214 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_213 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_212 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X4 FILL_211 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X4 FILL_210 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_209 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X4 FILL_208 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_207 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X8 FILL_206 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_205 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_204 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X8 FILL_203 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X8 FILL_202 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_201 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_200 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_199 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_198 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_197 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X4 FILL_196 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_195 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_194 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X4 FILL_193 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_192 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X4 FILL_191 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X8 FILL_190 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X32 FILL_189 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X4 FILL_188 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X4 FILL_187 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_186 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_185 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_184 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_183 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_182 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_181 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_180 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_179 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_178 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_177 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X4 FILL_176 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_175 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X4 FILL_174 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_173 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_172 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X8 FILL_171 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X8 FILL_170 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_169 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_168 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_167 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_166 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_165 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X16 FILL_164 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_163 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_162 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X4 FILL_161 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_160 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_159 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X8 FILL_158 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_157 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_156 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_155 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_154 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_153 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_152 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_151 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_150 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_149 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_148 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_147 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_146 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X4 FILL_145 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_144 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_143 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_142 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_141 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X4 FILL_140 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X16 FILL_139 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_138 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_137 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_136 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_135 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_134 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_133 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X4 FILL_132 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_131 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_130 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_129 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_128 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_127 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X4 FILL_126 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_125 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X4 FILL_124 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X4 FILL_123 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X8 FILL_122 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_121 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X4 FILL_120 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X8 FILL_119 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_118 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_117 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X4 FILL_116 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_115 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_114 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X4 FILL_113 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X4 FILL_112 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X8 FILL_111 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X32 FILL_110 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_109 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_108 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X4 FILL_107 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_106 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_105 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_104 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X4 FILL_103 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_102 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_101 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_100 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_99 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_98 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_97 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_96 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_95 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X4 FILL_94 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X16 FILL_93 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_92 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_91 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X4 FILL_90 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_89 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_88 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_87 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_86 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X4 FILL_85 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_84 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_83 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_82 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_81 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X4 FILL_80 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X8 FILL_79 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X16 FILL_78 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_77 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_76 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_75 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_74 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_73 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_72 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_71 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_70 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_69 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_68 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_67 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_66 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_65 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X4 FILL_64 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X8 FILL_63 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X16 FILL_62 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_61 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X4 FILL_60 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_59 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_58 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X4 FILL_57 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_56 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X4 FILL_55 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_54 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_53 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_52 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_51 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_50 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_49 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_48 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_47 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_46 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_45 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_44 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_43 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X4 FILL_42 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X4 FILL_41 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_40 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_39 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_38 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_37 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_36 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_35 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_34 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_33 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X4 FILL_32 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X32 FILL_31 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_30 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_29 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_28 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X8 FILL_27 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X4 FILL_26 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_25 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X4 FILL_24 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_23 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_22 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_21 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X4 FILL_20 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_19 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_18 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X4 FILL_17 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_16 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_15 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X4 FILL_14 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_13 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X8 FILL_12 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_11 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_10 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_9 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X4 FILL_8 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_7 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_6 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_5 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_4 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X2 FILL_3 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X4 FILL_2 (
	.VDD(VDD), 
	.VSS(VSS) );
   FILLCELL_X32 FILL_1 (
	.VDD(VDD), 
	.VSS(VSS) );
endmodule

