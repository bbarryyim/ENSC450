FLIP FLOP: Group 14 

* Technology Dependent design rules/parameters
.include /ensc/fac1/fcampi/esil/hspice/cmosp18/rules.inc

* Transistor models 
.protect
.LIB `/ensc/fac1/fcampi/esil/hspice/cmosp18/log018.l' TT  $ typical process corner.
.unprotect

* Supply Sources
.param pwr=1.2 
.temp  25
Vvdd  vdd  0 dc pwr
Vvdds vdds 0 dc pwr
Vgnd  gnd  0 dc 0
Vgnds gnds 0 dc 0

* Subcircuits
.subckt INV a z vdd gnd vdds gnds Wn=Wm#
Xpmos vdd a z vdds pt_st w=2*Wn
Xnmos gnd a z gnds nt_st w=Wn
.ends

.subckt TRANSGATE d g notg s vdds gnds Wn=Wm#  
Xnmos d g    s gnds nt_st w=Wn
Xpmos d notg s vdds pt_st wn=2*Wn
.ends

.subckt DLATCH d ck nck a notqm vdd gnd vdds gnds Wn=Wm#
Xtransgate1 d ck  nck a vdds gnds TRANSGATE Wn=Wm#
Xinv1 a     notqm vdd gnd vdds gnds INV Wn=Wm#
Xinv2 notqm b     vdd gnd vdds gnds INV Wn=Wm#
Xtransgate2 b nck ck  a vdds gnds TRANSGATE Wn=Wm#
.ends

* Logic 
.param Wn=Wm#
Xinvclk clk nclk vdd gnd vdds gnds INV Wn=Wm#
Xdlatch1 d    nclk clk  q     notq vdd gnd vdds gnds DLATCH Wn=Wm#
Xdlatch2 notq clk  nclk notq1 q1   vdd gnd vdds gnds DLATCH Wn=Wm#


Cload q1 0 20f

* Input Stimuli (Step response)
VD  	d  0 PWL(0n 0 0.7ns 0 0.8ns pwr 3.1ns pwr 3.2ns 0)
Vclk  clk  0 PWL(0n 0 0.4ns 0 0.5ns pwr 0.9ns pwr 1.0ns 0 1.4ns 0 1.5ns pwr 1.9ns pwr 2.0ns 0 2.4ns 0 2.5ns pwr 2.9ns pwr 3.0ns 0 3.4ns 0 3.5ns pwr 3.9ns pwr 4.0ns 0 4.4ns 0 4.5ns pwr 4.9ns pwr 5.0ns 0)

* Simulation Parameters ************************
*.tran 0.01ps 5.0ns START=0 

.tran 0.01ps 5.0ns START=0 sweep Wn START=Wm# STOP=300*Wm# STEP=50*Wm#

.option post
.meas tran tpd_in01      trig v(D) val='pwr*0.5' cross=1
+                        targ v(Q) val='pwr*0.5' cross=1 
.meas tran ttr           trig v(Q) val='pwr*0.8' fall=1
+                        targ v(Q) val='pwr*0.2' fall=1
.meas tran leak_pow_in1  avg power FROM=12ns TO=14ns
.meas tran leak_pow_in0  avg power FROM= 6ns TO= 8ns
.meas tran dyn_pow       avg power FROM= 9ns TO=10ns

************************************************

.end
  
